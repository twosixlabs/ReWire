module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [16:0] __in0,
  output logic [14:0] __out0);
  logic [90:0] zll_pure_dispatch7_in;
  logic [142:0] zll_pure_dispatch7_out;
  logic [90:0] zll_pure_dispatch8_in;
  logic [86:0] zll_main_reset10_in;
  logic [86:0] zll_main_putins5_in;
  logic [69:0] zll_main_putins5_out;
  logic [69:0] zll_main_loop226_in;
  logic [142:0] zll_main_loop226_out;
  logic [142:0] zll_main_reset39_in;
  logic [142:0] zll_main_reset30_in;
  logic [69:0] zll_main_reset32_in;
  logic [69:0] main_getpc_in;
  logic [75:0] main_getpc_out;
  logic [75:0] zll_main_loop135_in;
  logic [69:0] zll_main_loop135_out;
  logic [69:0] zll_main_loop226_inR1;
  logic [142:0] zll_main_loop226_outR1;
  logic [142:0] zll_main_reset46_in;
  logic [142:0] zll_main_reset35_in;
  logic [69:0] zll_main_reset34_in;
  logic [69:0] main_getout_in;
  logic [84:0] main_getout_out;
  logic [84:0] zll_main_loop197_in;
  logic [142:0] zll_main_loop197_out;
  logic [142:0] zll_main_reset44_in;
  logic [142:0] zll_main_reset26_in;
  logic [84:0] zll_main_reset17_in;
  logic [90:0] zll_pure_dispatch4_in;
  logic [86:0] zll_main_loop39_in;
  logic [86:0] zll_main_putins5_inR1;
  logic [69:0] zll_main_putins5_outR1;
  logic [69:0] zll_main_loop226_inR2;
  logic [142:0] zll_main_loop226_outR2;
  logic [142:0] zll_main_loop52_in;
  logic [142:0] zll_main_loop100_in;
  logic [69:0] zll_main_loop180_in;
  logic [69:0] main_incrpc_in;
  logic [69:0] main_incrpc_out;
  logic [69:0] zll_main_loop226_inR3;
  logic [142:0] zll_main_loop226_outR3;
  logic [142:0] zll_main_loop68_in;
  logic [142:0] zll_main_loop216_in;
  logic [69:0] zll_main_loop188_in;
  logic [69:0] main_getpc_inR1;
  logic [75:0] main_getpc_outR1;
  logic [75:0] zll_main_loop135_inR1;
  logic [69:0] zll_main_loop135_outR1;
  logic [69:0] zll_main_loop226_inR4;
  logic [142:0] zll_main_loop226_outR4;
  logic [142:0] zll_main_loop51_in;
  logic [142:0] zll_main_loop117_in;
  logic [69:0] zll_main_loop23_in;
  logic [69:0] main_getout_inR1;
  logic [84:0] main_getout_outR1;
  logic [84:0] zll_main_loop197_inR1;
  logic [142:0] zll_main_loop197_outR1;
  logic [142:0] zll_main_loop43_in;
  logic [142:0] zll_main_loop53_in;
  logic [84:0] zll_main_loop206_in;
  logic [90:0] zll_pure_dispatch7_inR1;
  logic [142:0] zll_pure_dispatch7_outR1;
  logic [90:0] zll_pure_dispatch7_inR2;
  logic [142:0] zll_pure_dispatch7_outR2;
  logic [90:0] zll_pure_dispatch3_in;
  logic [86:0] zll_main_loop132_in;
  logic [86:0] zll_main_putins5_inR2;
  logic [69:0] zll_main_putins5_outR2;
  logic [69:0] zll_main_loop226_inR5;
  logic [142:0] zll_main_loop226_outR5;
  logic [142:0] zll_main_loop190_in;
  logic [142:0] zll_main_loop107_in;
  logic [69:0] zll_main_loop159_in;
  logic [69:0] main_getdatain_in;
  logic [69:0] main_getins_in;
  logic [86:0] main_getins_out;
  logic [86:0] zll_main_getdatain1_in;
  logic [86:0] zll_main_getdatain_in;
  logic [16:0] zll_main_datain2_in;
  logic [16:0] zll_main_datain_in;
  logic [77:0] zll_main_loop16_in;
  logic [77:0] main_putreg_in;
  logic [89:0] zll_main_putreg15_in;
  logic [69:0] zll_main_putreg15_out;
  logic [69:0] zll_main_loop226_inR6;
  logic [142:0] zll_main_loop226_outR6;
  logic [142:0] zll_main_loop222_in;
  logic [142:0] zll_main_loop222_out;
  logic [90:0] zll_pure_dispatch6_in;
  logic [86:0] zll_main_loop155_in;
  logic [86:0] zll_main_putins5_inR3;
  logic [69:0] zll_main_putins5_outR3;
  logic [69:0] zll_main_loop226_inR7;
  logic [142:0] zll_main_loop226_outR7;
  logic [142:0] zll_main_loop141_in;
  logic [142:0] zll_main_loop6_in;
  logic [69:0] zll_main_loop211_in;
  logic [69:0] main_incrpc_inR1;
  logic [69:0] main_incrpc_outR1;
  logic [69:0] zll_main_loop226_inR8;
  logic [142:0] zll_main_loop226_outR8;
  logic [142:0] zll_main_loop31_in;
  logic [142:0] zll_main_loop214_in;
  logic [69:0] zll_main_loop179_in;
  logic [69:0] main_getpc_inR2;
  logic [75:0] main_getpc_outR2;
  logic [75:0] zll_main_loop135_inR2;
  logic [69:0] zll_main_loop135_outR2;
  logic [69:0] zll_main_loop226_inR9;
  logic [142:0] zll_main_loop226_outR9;
  logic [142:0] zll_main_loop213_in;
  logic [142:0] zll_main_loop120_in;
  logic [69:0] zll_main_loop158_in;
  logic [69:0] main_getout_inR2;
  logic [84:0] main_getout_outR2;
  logic [84:0] zll_main_loop197_inR2;
  logic [142:0] zll_main_loop197_outR2;
  logic [142:0] zll_main_loop119_in;
  logic [142:0] zll_main_loop47_in;
  logic [84:0] zll_main_loop87_in;
  logic [90:0] zll_pure_dispatch7_inR3;
  logic [142:0] zll_pure_dispatch7_outR3;
  logic [90:0] zll_pure_dispatch7_inR4;
  logic [142:0] zll_pure_dispatch7_outR4;
  logic [0:0] __continue;
  logic [52:0] __padding;
  logic [3:0] __resumption_tag;
  logic [69:0] __st0;
  logic [3:0] __resumption_tag_next;
  logic [69:0] __st0_next;
  assign zll_pure_dispatch7_in = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch7  inst (zll_pure_dispatch7_in[90:74], zll_pure_dispatch7_in[69:0], zll_pure_dispatch7_out);
  assign zll_pure_dispatch8_in = {__in0, {__resumption_tag, __st0}};
  assign zll_main_reset10_in = {zll_pure_dispatch8_in[90:74], zll_pure_dispatch8_in[69:0]};
  assign zll_main_putins5_in = {zll_main_reset10_in[86:70], zll_main_reset10_in[69:0]};
  ZLL_Main_putIns5  instR1 (zll_main_putins5_in[86:70], zll_main_putins5_in[69:0], zll_main_putins5_out);
  assign zll_main_loop226_in = zll_main_putins5_out;
  ZLL_Main_loop226  instR2 (zll_main_loop226_in[69:0], zll_main_loop226_out);
  assign zll_main_reset39_in = zll_main_loop226_out;
  assign zll_main_reset30_in = zll_main_reset39_in[142:0];
  assign zll_main_reset32_in = zll_main_reset30_in[69:0];
  assign main_getpc_in = zll_main_reset32_in[69:0];
  Main_getPC  instR3 (main_getpc_in[69:0], main_getpc_out);
  assign zll_main_loop135_in = main_getpc_out;
  ZLL_Main_loop135  instR4 (zll_main_loop135_in[75:0], zll_main_loop135_out);
  assign zll_main_loop226_inR1 = zll_main_loop135_out;
  ZLL_Main_loop226  instR5 (zll_main_loop226_inR1[69:0], zll_main_loop226_outR1);
  assign zll_main_reset46_in = zll_main_loop226_outR1;
  assign zll_main_reset35_in = zll_main_reset46_in[142:0];
  assign zll_main_reset34_in = zll_main_reset35_in[69:0];
  assign main_getout_in = zll_main_reset34_in[69:0];
  Main_getOut  instR6 (main_getout_in[69:0], main_getout_out);
  assign zll_main_loop197_in = main_getout_out;
  ZLL_Main_loop197  instR7 (zll_main_loop197_in[84:0], zll_main_loop197_out);
  assign zll_main_reset44_in = zll_main_loop197_out;
  assign zll_main_reset26_in = zll_main_reset44_in[142:0];
  assign zll_main_reset17_in = {zll_main_reset26_in[84:70], zll_main_reset26_in[69:0]};
  assign zll_pure_dispatch4_in = {__in0, {__resumption_tag, __st0}};
  assign zll_main_loop39_in = {zll_pure_dispatch4_in[90:74], zll_pure_dispatch4_in[69:0]};
  assign zll_main_putins5_inR1 = {zll_main_loop39_in[86:70], zll_main_loop39_in[69:0]};
  ZLL_Main_putIns5  instR8 (zll_main_putins5_inR1[86:70], zll_main_putins5_inR1[69:0], zll_main_putins5_outR1);
  assign zll_main_loop226_inR2 = zll_main_putins5_outR1;
  ZLL_Main_loop226  instR9 (zll_main_loop226_inR2[69:0], zll_main_loop226_outR2);
  assign zll_main_loop52_in = zll_main_loop226_outR2;
  assign zll_main_loop100_in = zll_main_loop52_in[142:0];
  assign zll_main_loop180_in = zll_main_loop100_in[69:0];
  assign main_incrpc_in = zll_main_loop180_in[69:0];
  Main_incrPC  instR10 (main_incrpc_in[69:0], main_incrpc_out);
  assign zll_main_loop226_inR3 = main_incrpc_out;
  ZLL_Main_loop226  instR11 (zll_main_loop226_inR3[69:0], zll_main_loop226_outR3);
  assign zll_main_loop68_in = zll_main_loop226_outR3;
  assign zll_main_loop216_in = zll_main_loop68_in[142:0];
  assign zll_main_loop188_in = zll_main_loop216_in[69:0];
  assign main_getpc_inR1 = zll_main_loop188_in[69:0];
  Main_getPC  instR12 (main_getpc_inR1[69:0], main_getpc_outR1);
  assign zll_main_loop135_inR1 = main_getpc_outR1;
  ZLL_Main_loop135  instR13 (zll_main_loop135_inR1[75:0], zll_main_loop135_outR1);
  assign zll_main_loop226_inR4 = zll_main_loop135_outR1;
  ZLL_Main_loop226  instR14 (zll_main_loop226_inR4[69:0], zll_main_loop226_outR4);
  assign zll_main_loop51_in = zll_main_loop226_outR4;
  assign zll_main_loop117_in = zll_main_loop51_in[142:0];
  assign zll_main_loop23_in = zll_main_loop117_in[69:0];
  assign main_getout_inR1 = zll_main_loop23_in[69:0];
  Main_getOut  instR15 (main_getout_inR1[69:0], main_getout_outR1);
  assign zll_main_loop197_inR1 = main_getout_outR1;
  ZLL_Main_loop197  instR16 (zll_main_loop197_inR1[84:0], zll_main_loop197_outR1);
  assign zll_main_loop43_in = zll_main_loop197_outR1;
  assign zll_main_loop53_in = zll_main_loop43_in[142:0];
  assign zll_main_loop206_in = {zll_main_loop53_in[84:70], zll_main_loop53_in[69:0]};
  assign zll_pure_dispatch7_inR1 = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch7  instR17 (zll_pure_dispatch7_inR1[90:74], zll_pure_dispatch7_inR1[69:0], zll_pure_dispatch7_outR1);
  assign zll_pure_dispatch7_inR2 = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch7  instR18 (zll_pure_dispatch7_inR2[90:74], zll_pure_dispatch7_inR2[69:0], zll_pure_dispatch7_outR2);
  assign zll_pure_dispatch3_in = {__in0, {__resumption_tag, __st0}};
  assign zll_main_loop132_in = {zll_pure_dispatch3_in[90:74], zll_pure_dispatch3_in[69:0]};
  assign zll_main_putins5_inR2 = {zll_main_loop132_in[86:70], zll_main_loop132_in[69:0]};
  ZLL_Main_putIns5  instR19 (zll_main_putins5_inR2[86:70], zll_main_putins5_inR2[69:0], zll_main_putins5_outR2);
  assign zll_main_loop226_inR5 = zll_main_putins5_outR2;
  ZLL_Main_loop226  instR20 (zll_main_loop226_inR5[69:0], zll_main_loop226_outR5);
  assign zll_main_loop190_in = zll_main_loop226_outR5;
  assign zll_main_loop107_in = zll_main_loop190_in[142:0];
  assign zll_main_loop159_in = zll_main_loop107_in[69:0];
  assign main_getdatain_in = zll_main_loop159_in[69:0];
  assign main_getins_in = main_getdatain_in[69:0];
  Main_getIns  instR21 (main_getins_in[69:0], main_getins_out);
  assign zll_main_getdatain1_in = main_getins_out;
  assign zll_main_getdatain_in = zll_main_getdatain1_in[86:0];
  assign zll_main_datain2_in = zll_main_getdatain_in[86:70];
  assign zll_main_datain_in = zll_main_datain2_in[16:0];
  assign zll_main_loop16_in = {zll_main_datain_in[7:0], zll_main_getdatain_in[69:0]};
  assign main_putreg_in = zll_main_loop16_in[77:0];
  assign zll_main_putreg15_in = {main_putreg_in[77:70], 4'h0, main_putreg_in[77:70], main_putreg_in[69:0]};
  ZLL_Main_putReg15  instR22 (zll_main_putreg15_in[89:82], zll_main_putreg15_in[81:80], zll_main_putreg15_in[79:70], zll_main_putreg15_in[69:0], zll_main_putreg15_out);
  assign zll_main_loop226_inR6 = zll_main_putreg15_out;
  ZLL_Main_loop226  instR23 (zll_main_loop226_inR6[69:0], zll_main_loop226_outR6);
  assign zll_main_loop222_in = zll_main_loop226_outR6;
  ZLL_Main_loop222  instR24 (zll_main_loop222_in[142:0], zll_main_loop222_out);
  assign zll_pure_dispatch6_in = {__in0, {__resumption_tag, __st0}};
  assign zll_main_loop155_in = {zll_pure_dispatch6_in[90:74], zll_pure_dispatch6_in[69:0]};
  assign zll_main_putins5_inR3 = {zll_main_loop155_in[86:70], zll_main_loop155_in[69:0]};
  ZLL_Main_putIns5  instR25 (zll_main_putins5_inR3[86:70], zll_main_putins5_inR3[69:0], zll_main_putins5_outR3);
  assign zll_main_loop226_inR7 = zll_main_putins5_outR3;
  ZLL_Main_loop226  instR26 (zll_main_loop226_inR7[69:0], zll_main_loop226_outR7);
  assign zll_main_loop141_in = zll_main_loop226_outR7;
  assign zll_main_loop6_in = zll_main_loop141_in[142:0];
  assign zll_main_loop211_in = zll_main_loop6_in[69:0];
  assign main_incrpc_inR1 = zll_main_loop211_in[69:0];
  Main_incrPC  instR27 (main_incrpc_inR1[69:0], main_incrpc_outR1);
  assign zll_main_loop226_inR8 = main_incrpc_outR1;
  ZLL_Main_loop226  instR28 (zll_main_loop226_inR8[69:0], zll_main_loop226_outR8);
  assign zll_main_loop31_in = zll_main_loop226_outR8;
  assign zll_main_loop214_in = zll_main_loop31_in[142:0];
  assign zll_main_loop179_in = zll_main_loop214_in[69:0];
  assign main_getpc_inR2 = zll_main_loop179_in[69:0];
  Main_getPC  instR29 (main_getpc_inR2[69:0], main_getpc_outR2);
  assign zll_main_loop135_inR2 = main_getpc_outR2;
  ZLL_Main_loop135  instR30 (zll_main_loop135_inR2[75:0], zll_main_loop135_outR2);
  assign zll_main_loop226_inR9 = zll_main_loop135_outR2;
  ZLL_Main_loop226  instR31 (zll_main_loop226_inR9[69:0], zll_main_loop226_outR9);
  assign zll_main_loop213_in = zll_main_loop226_outR9;
  assign zll_main_loop120_in = zll_main_loop213_in[142:0];
  assign zll_main_loop158_in = zll_main_loop120_in[69:0];
  assign main_getout_inR2 = zll_main_loop158_in[69:0];
  Main_getOut  instR32 (main_getout_inR2[69:0], main_getout_outR2);
  assign zll_main_loop197_inR2 = main_getout_outR2;
  ZLL_Main_loop197  instR33 (zll_main_loop197_inR2[84:0], zll_main_loop197_outR2);
  assign zll_main_loop119_in = zll_main_loop197_outR2;
  assign zll_main_loop47_in = zll_main_loop119_in[142:0];
  assign zll_main_loop87_in = {zll_main_loop47_in[84:70], zll_main_loop47_in[69:0]};
  assign zll_pure_dispatch7_inR3 = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch7  instR34 (zll_pure_dispatch7_inR3[90:74], zll_pure_dispatch7_inR3[69:0], zll_pure_dispatch7_outR3);
  assign zll_pure_dispatch7_inR4 = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch7  instR35 (zll_pure_dispatch7_inR4[90:74], zll_pure_dispatch7_inR4[69:0], zll_pure_dispatch7_outR4);
  assign {__continue, __padding, __out0, __resumption_tag_next, __st0_next} = (zll_pure_dispatch7_inR4[73:70] == 4'h1) ? zll_pure_dispatch7_outR4 : ((zll_pure_dispatch7_inR3[73:70] == 4'h2) ? zll_pure_dispatch7_outR3 : ((zll_pure_dispatch6_in[73:70] == 4'h3) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop87_in[84:70], 4'h4, zll_main_loop87_in[69:0]} : ((zll_pure_dispatch3_in[73:70] == 4'h4) ? zll_main_loop222_out : ((zll_pure_dispatch7_inR2[73:70] == 4'h5) ? zll_pure_dispatch7_outR2 : ((zll_pure_dispatch7_inR1[73:70] == 4'h6) ? zll_pure_dispatch7_outR1 : ((zll_pure_dispatch4_in[73:70] == 4'h7) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop206_in[84:70], 4'h0, zll_main_loop206_in[69:0]} : ((zll_pure_dispatch8_in[73:70] == 4'h8) ? {{1'h1, {6'h35{1'h0}}}, zll_main_reset17_in[84:70], 4'h1, zll_main_reset17_in[69:0]} : zll_pure_dispatch7_out)))))));
  initial {__resumption_tag, __st0} <= {1'h1, {7'h49{1'h0}}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      {__resumption_tag, __st0} <= {1'h1, {7'h49{1'h0}}};
    end else begin
      {__resumption_tag, __st0} <= {__resumption_tag_next, __st0_next};
    end
  end
endmodule

module ZLL_Main_loop226 (input logic [69:0] arg0,
  output logic [142:0] res);
  assign res = {{2'h1, {7'h47{1'h0}}}, arg0};
endmodule

module ZLL_Main_loop222 (input logic [142:0] arg0,
  output logic [142:0] res);
  logic [142:0] zll_main_reset42_in;
  logic [69:0] main_loop_in;
  logic [69:0] main_getinstr_in;
  logic [69:0] main_getins_in;
  logic [86:0] main_getins_out;
  logic [86:0] zll_main_getinstr1_in;
  logic [86:0] zll_main_getinstr2_in;
  logic [16:0] zll_main_instrin2_in;
  logic [16:0] zll_main_instrin1_in;
  logic [78:0] zll_main_loop113_in;
  logic [78:0] zll_main_loop136_in;
  logic [142:0] zll_main_loop59_in;
  logic [142:0] zll_main_loop173_in;
  logic [78:0] zll_main_loop171_in;
  logic [139:0] zll_main_loop124_in;
  logic [139:0] zll_main_loop218_in;
  logic [151:0] zll_main_loop143_in;
  logic [151:0] zll_main_loop154_in;
  logic [148:0] zll_main_loop_in;
  logic [78:0] zll_main_loop7_in;
  logic [75:0] zll_main_loop127_in;
  logic [75:0] zll_main_loop27_in;
  logic [69:0] main_getreg1_in;
  logic [77:0] main_getreg1_out;
  logic [83:0] zll_main_loop177_in;
  logic [83:0] zll_main_bnz_in;
  logic [15:0] binop_in;
  logic [84:0] zll_main_bnz1_in;
  logic [15:0] binop_inR1;
  logic [76:0] zll_main_bnz3_in;
  logic [76:0] zll_main_bnz5_in;
  logic [75:0] zll_main_bnz4_in;
  logic [75:0] zll_main_putpc12_in;
  logic [69:0] zll_main_putpc12_out;
  logic [70:0] zll_main_nand8_in;
  logic [69:0] main_incrpc_in;
  logic [69:0] main_incrpc_out;
  logic [69:0] zll_main_loop226_in;
  logic [142:0] zll_main_loop226_out;
  logic [142:0] zll_main_loop215_in;
  logic [142:0] zll_main_loop94_in;
  logic [69:0] zll_main_loop194_in;
  logic [69:0] main_getpc_in;
  logic [75:0] main_getpc_out;
  logic [75:0] zll_main_loop135_in;
  logic [69:0] zll_main_loop135_out;
  logic [69:0] zll_main_loop226_inR1;
  logic [142:0] zll_main_loop226_outR1;
  logic [142:0] zll_main_loop202_in;
  logic [142:0] zll_main_loop170_in;
  logic [69:0] zll_main_loop21_in;
  logic [69:0] main_getout_in;
  logic [84:0] main_getout_out;
  logic [84:0] zll_main_loop197_in;
  logic [142:0] zll_main_loop197_out;
  logic [142:0] zll_main_loop61_in;
  logic [142:0] zll_main_loop164_in;
  logic [84:0] zll_main_loop20_in;
  logic [78:0] zll_main_loop178_in;
  logic [75:0] zll_main_loop205_in;
  logic [75:0] zll_main_loop28_in;
  logic [75:0] zll_main_loop174_in;
  logic [75:0] zll_main_loop203_in;
  logic [71:0] main_getreg_in;
  logic [77:0] main_getreg_out;
  logic [81:0] zll_main_loop199_in;
  logic [81:0] zll_main_loop3_in;
  logic [81:0] zll_main_loop92_in;
  logic [81:0] zll_main_nand1_in;
  logic [71:0] main_getreg_inR1;
  logic [77:0] main_getreg_outR1;
  logic [87:0] zll_main_nand4_in;
  logic [87:0] zll_main_nand7_in;
  logic [87:0] zll_main_nand2_in;
  logic [87:0] zll_main_nand6_in;
  logic [15:0] binop_inR2;
  logic [7:0] unop_in;
  logic [79:0] main_putreg1_in;
  logic [89:0] zll_main_putreg15_in;
  logic [69:0] zll_main_putreg15_out;
  logic [69:0] main_incrpc_inR1;
  logic [69:0] main_incrpc_outR1;
  logic [69:0] zll_main_loop226_inR2;
  logic [142:0] zll_main_loop226_outR2;
  logic [142:0] zll_main_loop187_in;
  logic [142:0] zll_main_loop85_in;
  logic [69:0] zll_main_loop191_in;
  logic [69:0] main_getpc_inR1;
  logic [75:0] main_getpc_outR1;
  logic [75:0] zll_main_loop135_inR1;
  logic [69:0] zll_main_loop135_outR1;
  logic [69:0] zll_main_loop226_inR3;
  logic [142:0] zll_main_loop226_outR3;
  logic [142:0] zll_main_loop35_in;
  logic [142:0] zll_main_loop168_in;
  logic [69:0] zll_main_loop34_in;
  logic [69:0] main_getout_inR1;
  logic [84:0] main_getout_outR1;
  logic [84:0] zll_main_loop197_inR1;
  logic [142:0] zll_main_loop197_outR1;
  logic [142:0] zll_main_loop142_in;
  logic [142:0] zll_main_loop224_in;
  logic [84:0] zll_main_loop223_in;
  logic [78:0] zll_main_loop77_in;
  logic [75:0] zll_main_loop70_in;
  logic [75:0] zll_main_loop76_in;
  logic [69:0] main_getreg1_inR1;
  logic [77:0] main_getreg1_outR1;
  logic [83:0] zll_main_loop131_in;
  logic [83:0] zll_main_st9_in;
  logic [75:0] zll_main_putaddrout4_in;
  logic [69:0] zll_main_putaddrout4_out;
  logic [77:0] zll_main_st5_in;
  logic [77:0] zll_main_putdataout_in;
  logic [69:0] main_getout_inR2;
  logic [84:0] main_getout_outR2;
  logic [92:0] zll_main_putdataout1_in;
  logic [92:0] zll_main_putdataout5_in;
  logic [22:0] zll_main_putdataout9_in;
  logic [22:0] zll_main_putdataout2_in;
  logic [22:0] zll_main_putdataout4_in;
  logic [22:0] zll_main_putdataout10_in;
  logic [84:0] zll_main_putout12_in;
  logic [69:0] zll_main_putout12_out;
  logic [69:0] main_putweout_in;
  logic [70:0] zll_main_putweout6_in;
  logic [69:0] zll_main_putweout6_out;
  logic [69:0] zll_main_loop226_inR4;
  logic [142:0] zll_main_loop226_outR4;
  logic [142:0] zll_main_loop55_in;
  logic [142:0] zll_main_loop129_in;
  logic [69:0] zll_main_loop137_in;
  logic [69:0] main_getout_inR3;
  logic [84:0] main_getout_outR3;
  logic [84:0] zll_main_loop197_inR2;
  logic [142:0] zll_main_loop197_outR2;
  logic [142:0] zll_main_loop79_in;
  logic [142:0] zll_main_loop169_in;
  logic [84:0] zll_main_loop115_in;
  logic [78:0] zll_main_loop126_in;
  logic [75:0] zll_main_loop209_in;
  logic [75:0] zll_main_loop118_in;
  logic [75:0] zll_main_putaddrout4_inR1;
  logic [69:0] zll_main_putaddrout4_outR1;
  logic [69:0] main_putweout1_in;
  logic [69:0] main_putweout1_out;
  logic [69:0] zll_main_loop226_inR5;
  logic [142:0] zll_main_loop226_outR5;
  logic [142:0] zll_main_loop17_in;
  logic [142:0] zll_main_loop88_in;
  logic [69:0] zll_main_loop54_in;
  logic [69:0] main_getout_inR4;
  logic [84:0] main_getout_outR4;
  logic [84:0] zll_main_loop197_inR3;
  logic [142:0] zll_main_loop197_outR3;
  logic [142:0] zll_main_loop74_in;
  logic [142:0] zll_main_loop106_in;
  logic [84:0] zll_main_loop184_in;
  logic [78:0] zll_main_loop208_in;
  logic [69:0] zll_main_loop8_in;
  logic [69:0] main_incrpc_inR2;
  logic [69:0] main_incrpc_outR2;
  logic [69:0] zll_main_loop226_inR6;
  logic [142:0] zll_main_loop226_outR6;
  logic [142:0] zll_main_loop219_in;
  logic [142:0] zll_main_loop97_in;
  logic [69:0] zll_main_loop56_in;
  logic [69:0] main_getpc_inR2;
  logic [75:0] main_getpc_outR2;
  logic [75:0] zll_main_loop135_inR2;
  logic [69:0] zll_main_loop135_outR2;
  logic [69:0] zll_main_loop226_inR7;
  logic [142:0] zll_main_loop226_outR7;
  logic [142:0] zll_main_loop36_in;
  logic [142:0] zll_main_loop96_in;
  logic [69:0] zll_main_loop176_in;
  logic [69:0] main_getout_inR5;
  logic [84:0] main_getout_outR5;
  logic [84:0] zll_main_loop197_inR4;
  logic [142:0] zll_main_loop197_outR4;
  logic [142:0] zll_main_loop189_in;
  logic [142:0] zll_main_loop210_in;
  logic [84:0] zll_main_loop1_in;
  assign zll_main_reset42_in = arg0;
  assign main_loop_in = zll_main_reset42_in[69:0];
  assign main_getinstr_in = main_loop_in[69:0];
  assign main_getins_in = main_getinstr_in[69:0];
  Main_getIns  inst (main_getins_in[69:0], main_getins_out);
  assign zll_main_getinstr1_in = main_getins_out;
  assign zll_main_getinstr2_in = zll_main_getinstr1_in[86:0];
  assign zll_main_instrin2_in = zll_main_getinstr2_in[86:70];
  assign zll_main_instrin1_in = zll_main_instrin2_in[16:0];
  assign zll_main_loop113_in = {zll_main_instrin1_in[16:8], zll_main_getinstr2_in[69:0]};
  assign zll_main_loop136_in = zll_main_loop113_in[78:0];
  assign zll_main_loop59_in = {{7'h40{1'h0}}, zll_main_loop136_in[78:70], zll_main_loop136_in[69:0]};
  assign zll_main_loop173_in = zll_main_loop59_in[142:0];
  assign zll_main_loop171_in = {zll_main_loop173_in[78:70], zll_main_loop173_in[69:0]};
  assign zll_main_loop124_in = {zll_main_loop171_in[69:0], zll_main_loop171_in[69:0]};
  assign zll_main_loop218_in = zll_main_loop124_in[139:0];
  assign zll_main_loop143_in = {zll_main_loop171_in[78:70], {3'h3, zll_main_loop218_in[139:70], zll_main_loop218_in[69:0]}};
  assign zll_main_loop154_in = {zll_main_loop143_in[151:143], zll_main_loop143_in[142:0]};
  assign zll_main_loop_in = {zll_main_loop154_in[151:143], zll_main_loop154_in[139:70], zll_main_loop154_in[69:0]};
  assign zll_main_loop7_in = {zll_main_loop_in[69:0], zll_main_loop_in[148:140]};
  assign zll_main_loop127_in = {zll_main_loop7_in[78:9], zll_main_loop7_in[5:0]};
  assign zll_main_loop27_in = {zll_main_loop127_in[5:0], zll_main_loop127_in[75:6]};
  assign main_getreg1_in = zll_main_loop27_in[69:0];
  Main_getReg1  instR1 (main_getreg1_in[69:0], main_getreg1_out);
  assign zll_main_loop177_in = {zll_main_loop27_in[75:70], main_getreg1_out};
  assign zll_main_bnz_in = {zll_main_loop177_in[83:78], zll_main_loop177_in[77:0]};
  assign binop_in = {zll_main_bnz_in[77:70], 8'h0};
  assign zll_main_bnz1_in = {zll_main_bnz_in[83:78], zll_main_bnz_in[77:70], binop_in[15:8] == binop_in[7:0], zll_main_bnz_in[69:0]};
  assign binop_inR1 = {zll_main_bnz1_in[78:71], 8'h0};
  assign zll_main_bnz3_in = {zll_main_bnz1_in[84:79], binop_inR1[15:8] == binop_inR1[7:0], zll_main_bnz1_in[69:0]};
  assign zll_main_bnz5_in = {zll_main_bnz3_in[69:0], zll_main_bnz3_in[76:71], zll_main_bnz3_in[70]};
  assign zll_main_bnz4_in = {zll_main_bnz5_in[76:7], zll_main_bnz5_in[6:1]};
  assign zll_main_putpc12_in = {zll_main_bnz4_in[5:0], zll_main_bnz4_in[75:6]};
  ZLL_Main_putPC12  instR2 (zll_main_putpc12_in[75:70], zll_main_putpc12_in[69:0], zll_main_putpc12_out);
  assign zll_main_nand8_in = {zll_main_bnz1_in[69:0], zll_main_bnz1_in[70]};
  assign main_incrpc_in = zll_main_nand8_in[70:1];
  Main_incrPC  instR3 (main_incrpc_in[69:0], main_incrpc_out);
  assign zll_main_loop226_in = (zll_main_nand8_in[0] == 1'h1) ? main_incrpc_out : zll_main_putpc12_out;
  ZLL_Main_loop226  instR4 (zll_main_loop226_in[69:0], zll_main_loop226_out);
  assign zll_main_loop215_in = zll_main_loop226_out;
  assign zll_main_loop94_in = zll_main_loop215_in[142:0];
  assign zll_main_loop194_in = zll_main_loop94_in[69:0];
  assign main_getpc_in = zll_main_loop194_in[69:0];
  Main_getPC  instR5 (main_getpc_in[69:0], main_getpc_out);
  assign zll_main_loop135_in = main_getpc_out;
  ZLL_Main_loop135  instR6 (zll_main_loop135_in[75:0], zll_main_loop135_out);
  assign zll_main_loop226_inR1 = zll_main_loop135_out;
  ZLL_Main_loop226  instR7 (zll_main_loop226_inR1[69:0], zll_main_loop226_outR1);
  assign zll_main_loop202_in = zll_main_loop226_outR1;
  assign zll_main_loop170_in = zll_main_loop202_in[142:0];
  assign zll_main_loop21_in = zll_main_loop170_in[69:0];
  assign main_getout_in = zll_main_loop21_in[69:0];
  Main_getOut  instR8 (main_getout_in[69:0], main_getout_out);
  assign zll_main_loop197_in = main_getout_out;
  ZLL_Main_loop197  instR9 (zll_main_loop197_in[84:0], zll_main_loop197_out);
  assign zll_main_loop61_in = zll_main_loop197_out;
  assign zll_main_loop164_in = zll_main_loop61_in[142:0];
  assign zll_main_loop20_in = {zll_main_loop164_in[84:70], zll_main_loop164_in[69:0]};
  assign zll_main_loop178_in = {zll_main_loop_in[69:0], zll_main_loop_in[148:140]};
  assign zll_main_loop205_in = {zll_main_loop178_in[78:9], zll_main_loop178_in[5:4], zll_main_loop178_in[3:2], zll_main_loop178_in[1:0]};
  assign zll_main_loop28_in = {zll_main_loop205_in[75:6], zll_main_loop205_in[3:2], zll_main_loop205_in[5:4], zll_main_loop205_in[1:0]};
  assign zll_main_loop174_in = {zll_main_loop28_in[3:2], zll_main_loop28_in[5:4], zll_main_loop28_in[1:0], zll_main_loop28_in[75:6]};
  assign zll_main_loop203_in = {zll_main_loop174_in[73:72], zll_main_loop174_in[75:74], zll_main_loop174_in[71:70], zll_main_loop174_in[69:0]};
  assign main_getreg_in = {zll_main_loop203_in[75:74], zll_main_loop203_in[69:0]};
  Main_getReg  instR10 (main_getreg_in[71:70], main_getreg_in[69:0], main_getreg_out);
  assign zll_main_loop199_in = {zll_main_loop203_in[73:72], zll_main_loop203_in[71:70], main_getreg_out};
  assign zll_main_loop3_in = {zll_main_loop199_in[81:80], zll_main_loop199_in[79:78], zll_main_loop199_in[77:0]};
  assign zll_main_loop92_in = {zll_main_loop3_in[79:78], zll_main_loop3_in[81:80], zll_main_loop3_in[77:70], zll_main_loop3_in[69:0]};
  assign zll_main_nand1_in = {zll_main_loop92_in[79:78], zll_main_loop92_in[81:80], zll_main_loop92_in[77:70], zll_main_loop92_in[69:0]};
  assign main_getreg_inR1 = {zll_main_nand1_in[79:78], zll_main_nand1_in[69:0]};
  Main_getReg  instR11 (main_getreg_inR1[71:70], main_getreg_inR1[69:0], main_getreg_outR1);
  assign zll_main_nand4_in = {zll_main_nand1_in[81:80], zll_main_nand1_in[77:70], main_getreg_outR1};
  assign zll_main_nand7_in = {zll_main_nand4_in[87:86], zll_main_nand4_in[85:78], zll_main_nand4_in[77:0]};
  assign zll_main_nand2_in = {zll_main_nand7_in[85:78], zll_main_nand7_in[87:86], zll_main_nand7_in[77:70], zll_main_nand7_in[69:0]};
  assign zll_main_nand6_in = {zll_main_nand2_in[79:78], zll_main_nand2_in[87:80], zll_main_nand2_in[77:70], zll_main_nand2_in[69:0]};
  assign binop_inR2 = {zll_main_nand6_in[85:78], zll_main_nand6_in[77:70]};
  assign unop_in = binop_inR2[15:8] & binop_inR2[7:0];
  assign main_putreg1_in = {zll_main_nand6_in[87:86], ~unop_in[7:0], zll_main_nand6_in[69:0]};
  assign zll_main_putreg15_in = {main_putreg1_in[77:70], main_putreg1_in[79:78], main_putreg1_in[79:78], main_putreg1_in[77:70], main_putreg1_in[69:0]};
  ZLL_Main_putReg15  instR12 (zll_main_putreg15_in[89:82], zll_main_putreg15_in[81:80], zll_main_putreg15_in[79:70], zll_main_putreg15_in[69:0], zll_main_putreg15_out);
  assign main_incrpc_inR1 = zll_main_putreg15_out;
  Main_incrPC  instR13 (main_incrpc_inR1[69:0], main_incrpc_outR1);
  assign zll_main_loop226_inR2 = main_incrpc_outR1;
  ZLL_Main_loop226  instR14 (zll_main_loop226_inR2[69:0], zll_main_loop226_outR2);
  assign zll_main_loop187_in = zll_main_loop226_outR2;
  assign zll_main_loop85_in = zll_main_loop187_in[142:0];
  assign zll_main_loop191_in = zll_main_loop85_in[69:0];
  assign main_getpc_inR1 = zll_main_loop191_in[69:0];
  Main_getPC  instR15 (main_getpc_inR1[69:0], main_getpc_outR1);
  assign zll_main_loop135_inR1 = main_getpc_outR1;
  ZLL_Main_loop135  instR16 (zll_main_loop135_inR1[75:0], zll_main_loop135_outR1);
  assign zll_main_loop226_inR3 = zll_main_loop135_outR1;
  ZLL_Main_loop226  instR17 (zll_main_loop226_inR3[69:0], zll_main_loop226_outR3);
  assign zll_main_loop35_in = zll_main_loop226_outR3;
  assign zll_main_loop168_in = zll_main_loop35_in[142:0];
  assign zll_main_loop34_in = zll_main_loop168_in[69:0];
  assign main_getout_inR1 = zll_main_loop34_in[69:0];
  Main_getOut  instR18 (main_getout_inR1[69:0], main_getout_outR1);
  assign zll_main_loop197_inR1 = main_getout_outR1;
  ZLL_Main_loop197  instR19 (zll_main_loop197_inR1[84:0], zll_main_loop197_outR1);
  assign zll_main_loop142_in = zll_main_loop197_outR1;
  assign zll_main_loop224_in = zll_main_loop142_in[142:0];
  assign zll_main_loop223_in = {zll_main_loop224_in[84:70], zll_main_loop224_in[69:0]};
  assign zll_main_loop77_in = {zll_main_loop_in[69:0], zll_main_loop_in[148:140]};
  assign zll_main_loop70_in = {zll_main_loop77_in[78:9], zll_main_loop77_in[5:0]};
  assign zll_main_loop76_in = {zll_main_loop70_in[5:0], zll_main_loop70_in[75:6]};
  assign main_getreg1_inR1 = zll_main_loop76_in[69:0];
  Main_getReg1  instR20 (main_getreg1_inR1[69:0], main_getreg1_outR1);
  assign zll_main_loop131_in = {zll_main_loop76_in[75:70], main_getreg1_outR1};
  assign zll_main_st9_in = {zll_main_loop131_in[83:78], zll_main_loop131_in[77:0]};
  assign zll_main_putaddrout4_in = {zll_main_st9_in[83:78], zll_main_st9_in[69:0]};
  ZLL_Main_putAddrOut4  instR21 (zll_main_putaddrout4_in[75:70], zll_main_putaddrout4_in[69:0], zll_main_putaddrout4_out);
  assign zll_main_st5_in = {zll_main_st9_in[77:70], zll_main_putaddrout4_out};
  assign zll_main_putdataout_in = {zll_main_st5_in[77:70], zll_main_st5_in[69:0]};
  assign main_getout_inR2 = zll_main_putdataout_in[69:0];
  Main_getOut  instR22 (main_getout_inR2[69:0], main_getout_outR2);
  assign zll_main_putdataout1_in = {zll_main_putdataout_in[77:70], main_getout_outR2};
  assign zll_main_putdataout5_in = {zll_main_putdataout1_in[92:85], zll_main_putdataout1_in[84:0]};
  assign zll_main_putdataout9_in = {zll_main_putdataout5_in[92:85], zll_main_putdataout5_in[84:70]};
  assign zll_main_putdataout2_in = {zll_main_putdataout9_in[22:15], zll_main_putdataout9_in[14:0]};
  assign zll_main_putdataout4_in = {zll_main_putdataout2_in[14], zll_main_putdataout2_in[22:15], zll_main_putdataout2_in[13:8], zll_main_putdataout2_in[7:0]};
  assign zll_main_putdataout10_in = {zll_main_putdataout4_in[13:8], zll_main_putdataout4_in[22], zll_main_putdataout4_in[21:14], zll_main_putdataout4_in[7:0]};
  assign zll_main_putout12_in = {{zll_main_putdataout10_in[16], zll_main_putdataout10_in[22:17], zll_main_putdataout10_in[15:8]}, zll_main_putdataout5_in[69:0]};
  ZLL_Main_putOut12  instR23 (zll_main_putout12_in[84:70], zll_main_putout12_in[69:0], zll_main_putout12_out);
  assign main_putweout_in = zll_main_putout12_out;
  assign zll_main_putweout6_in = {1'h1, main_putweout_in[69:0]};
  ZLL_Main_putWeOut6  instR24 (zll_main_putweout6_in[70], zll_main_putweout6_in[69:0], zll_main_putweout6_out);
  assign zll_main_loop226_inR4 = zll_main_putweout6_out;
  ZLL_Main_loop226  instR25 (zll_main_loop226_inR4[69:0], zll_main_loop226_outR4);
  assign zll_main_loop55_in = zll_main_loop226_outR4;
  assign zll_main_loop129_in = zll_main_loop55_in[142:0];
  assign zll_main_loop137_in = zll_main_loop129_in[69:0];
  assign main_getout_inR3 = zll_main_loop137_in[69:0];
  Main_getOut  instR26 (main_getout_inR3[69:0], main_getout_outR3);
  assign zll_main_loop197_inR2 = main_getout_outR3;
  ZLL_Main_loop197  instR27 (zll_main_loop197_inR2[84:0], zll_main_loop197_outR2);
  assign zll_main_loop79_in = zll_main_loop197_outR2;
  assign zll_main_loop169_in = zll_main_loop79_in[142:0];
  assign zll_main_loop115_in = {zll_main_loop169_in[84:70], zll_main_loop169_in[69:0]};
  assign zll_main_loop126_in = {zll_main_loop_in[69:0], zll_main_loop_in[148:140]};
  assign zll_main_loop209_in = {zll_main_loop126_in[78:9], zll_main_loop126_in[5:0]};
  assign zll_main_loop118_in = {zll_main_loop209_in[5:0], zll_main_loop209_in[75:6]};
  assign zll_main_putaddrout4_inR1 = {zll_main_loop118_in[75:70], zll_main_loop118_in[69:0]};
  ZLL_Main_putAddrOut4  instR28 (zll_main_putaddrout4_inR1[75:70], zll_main_putaddrout4_inR1[69:0], zll_main_putaddrout4_outR1);
  assign main_putweout1_in = zll_main_putaddrout4_outR1;
  Main_putWeOut1  instR29 (main_putweout1_in[69:0], main_putweout1_out);
  assign zll_main_loop226_inR5 = main_putweout1_out;
  ZLL_Main_loop226  instR30 (zll_main_loop226_inR5[69:0], zll_main_loop226_outR5);
  assign zll_main_loop17_in = zll_main_loop226_outR5;
  assign zll_main_loop88_in = zll_main_loop17_in[142:0];
  assign zll_main_loop54_in = zll_main_loop88_in[69:0];
  assign main_getout_inR4 = zll_main_loop54_in[69:0];
  Main_getOut  instR31 (main_getout_inR4[69:0], main_getout_outR4);
  assign zll_main_loop197_inR3 = main_getout_outR4;
  ZLL_Main_loop197  instR32 (zll_main_loop197_inR3[84:0], zll_main_loop197_outR3);
  assign zll_main_loop74_in = zll_main_loop197_outR3;
  assign zll_main_loop106_in = zll_main_loop74_in[142:0];
  assign zll_main_loop184_in = {zll_main_loop106_in[84:70], zll_main_loop106_in[69:0]};
  assign zll_main_loop208_in = {zll_main_loop_in[69:0], zll_main_loop_in[148:140]};
  assign zll_main_loop8_in = zll_main_loop208_in[78:9];
  assign main_incrpc_inR2 = zll_main_loop8_in[69:0];
  Main_incrPC  instR33 (main_incrpc_inR2[69:0], main_incrpc_outR2);
  assign zll_main_loop226_inR6 = main_incrpc_outR2;
  ZLL_Main_loop226  instR34 (zll_main_loop226_inR6[69:0], zll_main_loop226_outR6);
  assign zll_main_loop219_in = zll_main_loop226_outR6;
  assign zll_main_loop97_in = zll_main_loop219_in[142:0];
  assign zll_main_loop56_in = zll_main_loop97_in[69:0];
  assign main_getpc_inR2 = zll_main_loop56_in[69:0];
  Main_getPC  instR35 (main_getpc_inR2[69:0], main_getpc_outR2);
  assign zll_main_loop135_inR2 = main_getpc_outR2;
  ZLL_Main_loop135  instR36 (zll_main_loop135_inR2[75:0], zll_main_loop135_outR2);
  assign zll_main_loop226_inR7 = zll_main_loop135_outR2;
  ZLL_Main_loop226  instR37 (zll_main_loop226_inR7[69:0], zll_main_loop226_outR7);
  assign zll_main_loop36_in = zll_main_loop226_outR7;
  assign zll_main_loop96_in = zll_main_loop36_in[142:0];
  assign zll_main_loop176_in = zll_main_loop96_in[69:0];
  assign main_getout_inR5 = zll_main_loop176_in[69:0];
  Main_getOut  instR38 (main_getout_inR5[69:0], main_getout_outR5);
  assign zll_main_loop197_inR4 = main_getout_outR5;
  ZLL_Main_loop197  instR39 (zll_main_loop197_inR4[84:0], zll_main_loop197_outR4);
  assign zll_main_loop189_in = zll_main_loop197_outR4;
  assign zll_main_loop210_in = zll_main_loop189_in[142:0];
  assign zll_main_loop1_in = {zll_main_loop210_in[84:70], zll_main_loop210_in[69:0]};
  assign res = (zll_main_loop208_in[8:6] == 3'h0) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop1_in[84:70], 4'h6, zll_main_loop1_in[69:0]} : ((zll_main_loop126_in[8:6] == 3'h1) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop184_in[84:70], 4'h3, zll_main_loop184_in[69:0]} : ((zll_main_loop77_in[8:6] == 3'h2) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop115_in[84:70], 4'h7, zll_main_loop115_in[69:0]} : ((zll_main_loop178_in[8:6] == 3'h3) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop223_in[84:70], 4'h2, zll_main_loop223_in[69:0]} : {{1'h1, {6'h35{1'h0}}}, zll_main_loop20_in[84:70], 4'h5, zll_main_loop20_in[69:0]})));
endmodule

module ZLL_Main_putPC12 (input logic [5:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [145:0] zll_main_putpc10_in;
  logic [145:0] zll_main_putpc11_in;
  logic [75:0] zll_main_putpc13_in;
  logic [75:0] zll_main_putpc8_in;
  logic [75:0] zll_main_putpc2_in;
  logic [75:0] zll_main_putpc3_in;
  logic [75:0] zll_main_putpc_in;
  logic [69:0] zll_main_putpc14_in;
  assign zll_main_putpc10_in = {arg0, arg1, arg1};
  assign zll_main_putpc11_in = {zll_main_putpc10_in[145:140], zll_main_putpc10_in[139:0]};
  assign zll_main_putpc13_in = {zll_main_putpc11_in[145:140], zll_main_putpc11_in[139:70]};
  assign zll_main_putpc8_in = {zll_main_putpc13_in[75:70], zll_main_putpc13_in[69:0]};
  assign zll_main_putpc2_in = {zll_main_putpc8_in[69:62], zll_main_putpc8_in[75:70], zll_main_putpc8_in[61:54], zll_main_putpc8_in[53:46], zll_main_putpc8_in[45:38], zll_main_putpc8_in[37:32], zll_main_putpc8_in[31:15], zll_main_putpc8_in[14:0]};
  assign zll_main_putpc3_in = {zll_main_putpc2_in[61:54], zll_main_putpc2_in[75:68], zll_main_putpc2_in[67:62], zll_main_putpc2_in[53:46], zll_main_putpc2_in[45:38], zll_main_putpc2_in[37:32], zll_main_putpc2_in[31:15], zll_main_putpc2_in[14:0]};
  assign zll_main_putpc_in = {zll_main_putpc3_in[75:68], zll_main_putpc3_in[67:60], zll_main_putpc3_in[45:38], zll_main_putpc3_in[59:54], zll_main_putpc3_in[53:46], zll_main_putpc3_in[37:32], zll_main_putpc3_in[31:15], zll_main_putpc3_in[14:0]};
  assign zll_main_putpc14_in = {zll_main_putpc_in[75:68], zll_main_putpc_in[67:60], zll_main_putpc_in[59:52], zll_main_putpc_in[51:46], zll_main_putpc_in[45:38], zll_main_putpc_in[31:15], zll_main_putpc_in[14:0]};
  assign res = {zll_main_putpc14_in[61:54], zll_main_putpc14_in[69:62], zll_main_putpc14_in[39:32], zll_main_putpc14_in[53:46], zll_main_putpc14_in[45:40], zll_main_putpc14_in[31:15], zll_main_putpc14_in[14:0]};
endmodule

module ZLL_Main_putOut12 (input logic [14:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [154:0] zll_main_putout9_in;
  logic [154:0] zll_main_putout_in;
  logic [84:0] zll_main_putout5_in;
  logic [84:0] zll_main_putout7_in;
  logic [84:0] zll_main_putout14_in;
  logic [84:0] zll_main_putout11_in;
  logic [84:0] zll_main_putout8_in;
  assign zll_main_putout9_in = {arg0, arg1, arg1};
  assign zll_main_putout_in = {zll_main_putout9_in[154:140], zll_main_putout9_in[139:0]};
  assign zll_main_putout5_in = {zll_main_putout_in[154:140], zll_main_putout_in[139:70]};
  assign zll_main_putout7_in = {zll_main_putout5_in[84:70], zll_main_putout5_in[69:0]};
  assign zll_main_putout14_in = {zll_main_putout7_in[53:46], zll_main_putout7_in[84:70], zll_main_putout7_in[69:62], zll_main_putout7_in[61:54], zll_main_putout7_in[45:38], zll_main_putout7_in[37:32], zll_main_putout7_in[31:15], zll_main_putout7_in[14:0]};
  assign zll_main_putout11_in = {zll_main_putout14_in[45:38], zll_main_putout14_in[84:77], zll_main_putout14_in[76:62], zll_main_putout14_in[61:54], zll_main_putout14_in[53:46], zll_main_putout14_in[37:32], zll_main_putout14_in[31:15], zll_main_putout14_in[14:0]};
  assign zll_main_putout8_in = {zll_main_putout11_in[84:77], zll_main_putout11_in[76:69], zll_main_putout11_in[37:32], zll_main_putout11_in[68:54], zll_main_putout11_in[53:46], zll_main_putout11_in[45:38], zll_main_putout11_in[31:15], zll_main_putout11_in[14:0]};
  assign res = {zll_main_putout8_in[47:40], zll_main_putout8_in[39:32], zll_main_putout8_in[76:69], zll_main_putout8_in[84:77], zll_main_putout8_in[68:63], zll_main_putout8_in[31:15], zll_main_putout8_in[62:48]};
endmodule

module ZLL_Main_r17 (input logic [7:0] arg0,
  input logic [7:0] arg1,
  input logic [7:0] arg2,
  input logic [5:0] arg3,
  input logic [16:0] arg4,
  input logic [14:0] arg5,
  output logic [7:0] res);
  logic [53:0] zll_main_r07_in;
  logic [7:0] zll_main_r07_out;
  assign zll_main_r07_in = {arg0, arg2, arg3, arg4, arg5};
  ZLL_Main_r07  inst (zll_main_r07_in[53:46], zll_main_r07_in[45:38], zll_main_r07_in[37:32], zll_main_r07_in[31:15], zll_main_r07_in[14:0], zll_main_r07_out);
  assign res = zll_main_r07_out;
endmodule

module ZLL_Main_loop197 (input logic [84:0] arg0,
  output logic [142:0] res);
  logic [84:0] zll_main_loop175_in;
  assign zll_main_loop175_in = arg0;
  assign res = {{3'h1, {6'h37{1'h0}}}, zll_main_loop175_in[84:70], zll_main_loop175_in[69:0]};
endmodule

module ZLL_Main_r07 (input logic [7:0] arg0,
  input logic [7:0] arg1,
  input logic [5:0] arg2,
  input logic [16:0] arg3,
  input logic [14:0] arg4,
  output logic [7:0] res);
  logic [45:0] zll_main_r35_in;
  logic [7:0] zll_main_r35_out;
  assign zll_main_r35_in = {arg0, arg2, arg3, arg4};
  ZLL_Main_r35  inst (zll_main_r35_in[45:38], zll_main_r35_in[37:32], zll_main_r35_in[31:15], zll_main_r35_in[14:0], zll_main_r35_out);
  assign res = zll_main_r35_out;
endmodule

module ZLL_Main_r35 (input logic [7:0] arg0,
  input logic [5:0] arg1,
  input logic [16:0] arg2,
  input logic [14:0] arg3,
  output logic [7:0] res);
  logic [39:0] zll_main_r04_in;
  logic [22:0] zll_main_r27_in;
  assign zll_main_r04_in = {arg0, arg2, arg3};
  assign zll_main_r27_in = {zll_main_r04_in[39:32], zll_main_r04_in[14:0]};
  assign res = zll_main_r27_in[22:15];
endmodule

module Main_getReg1 (input logic [69:0] arg0,
  output logic [77:0] res);
  logic [73:0] zll_main_getreg13_in;
  logic [77:0] zll_main_getreg13_out;
  assign zll_main_getreg13_in = {4'h0, arg0};
  ZLL_Main_getReg13  inst (zll_main_getreg13_in[73:72], zll_main_getreg13_in[71:70], zll_main_getreg13_in[69:0], zll_main_getreg13_out);
  assign res = zll_main_getreg13_out;
endmodule

module Main_getReg (input logic [1:0] arg0,
  input logic [69:0] arg1,
  output logic [77:0] res);
  logic [73:0] zll_main_getreg13_in;
  logic [77:0] zll_main_getreg13_out;
  assign zll_main_getreg13_in = {arg0, arg0, arg1};
  ZLL_Main_getReg13  inst (zll_main_getreg13_in[73:72], zll_main_getreg13_in[71:70], zll_main_getreg13_in[69:0], zll_main_getreg13_out);
  assign res = zll_main_getreg13_out;
endmodule

module ZLL_Main_putWeOut6 (input logic [0:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [69:0] main_getout_in;
  logic [84:0] main_getout_out;
  logic [85:0] zll_main_putweout8_in;
  logic [85:0] zll_main_putweout1_in;
  logic [15:0] zll_main_putweout9_in;
  logic [15:0] zll_main_putweout7_in;
  logic [84:0] zll_main_putout12_in;
  logic [69:0] zll_main_putout12_out;
  assign main_getout_in = arg1;
  Main_getOut  inst (main_getout_in[69:0], main_getout_out);
  assign zll_main_putweout8_in = {arg0, main_getout_out};
  assign zll_main_putweout1_in = {zll_main_putweout8_in[85], zll_main_putweout8_in[84:0]};
  assign zll_main_putweout9_in = {zll_main_putweout1_in[85], zll_main_putweout1_in[84:70]};
  assign zll_main_putweout7_in = {zll_main_putweout9_in[15], zll_main_putweout9_in[14:0]};
  assign zll_main_putout12_in = {{zll_main_putweout7_in[15], zll_main_putweout7_in[13:8], zll_main_putweout7_in[7:0]}, zll_main_putweout1_in[69:0]};
  ZLL_Main_putOut12  instR1 (zll_main_putout12_in[84:70], zll_main_putout12_in[69:0], zll_main_putout12_out);
  assign res = zll_main_putout12_out;
endmodule

module Main_getIns (input logic [69:0] arg0,
  output logic [86:0] res);
  logic [139:0] zll_main_getins1_in;
  logic [139:0] zll_main_getins_in;
  logic [69:0] zll_main_inputs1_in;
  logic [69:0] zll_main_inputs5_in;
  logic [61:0] zll_main_inputs6_in;
  logic [53:0] zll_main_inputs2_in;
  logic [45:0] zll_main_inputs3_in;
  logic [37:0] zll_main_inputs4_in;
  logic [31:0] zll_main_inputs7_in;
  assign zll_main_getins1_in = {arg0, arg0};
  assign zll_main_getins_in = zll_main_getins1_in[139:0];
  assign zll_main_inputs1_in = zll_main_getins_in[139:70];
  assign zll_main_inputs5_in = zll_main_inputs1_in[69:0];
  assign zll_main_inputs6_in = {zll_main_inputs5_in[61:54], zll_main_inputs5_in[53:46], zll_main_inputs5_in[45:38], zll_main_inputs5_in[37:32], zll_main_inputs5_in[31:15], zll_main_inputs5_in[14:0]};
  assign zll_main_inputs2_in = {zll_main_inputs6_in[53:46], zll_main_inputs6_in[45:38], zll_main_inputs6_in[37:32], zll_main_inputs6_in[31:15], zll_main_inputs6_in[14:0]};
  assign zll_main_inputs3_in = {zll_main_inputs2_in[45:38], zll_main_inputs2_in[37:32], zll_main_inputs2_in[31:15], zll_main_inputs2_in[14:0]};
  assign zll_main_inputs4_in = {zll_main_inputs3_in[37:32], zll_main_inputs3_in[31:15], zll_main_inputs3_in[14:0]};
  assign zll_main_inputs7_in = {zll_main_inputs4_in[31:15], zll_main_inputs4_in[14:0]};
  assign res = {zll_main_inputs7_in[31:15], zll_main_getins_in[69:0]};
endmodule

module ZLL_Main_putAddrOut4 (input logic [5:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [69:0] main_getout_in;
  logic [84:0] main_getout_out;
  logic [90:0] zll_main_putaddrout7_in;
  logic [90:0] zll_main_putaddrout2_in;
  logic [20:0] zll_main_putaddrout6_in;
  logic [20:0] zll_main_putaddrout1_in;
  logic [84:0] zll_main_putout12_in;
  logic [69:0] zll_main_putout12_out;
  assign main_getout_in = arg1;
  Main_getOut  inst (main_getout_in[69:0], main_getout_out);
  assign zll_main_putaddrout7_in = {arg0, main_getout_out};
  assign zll_main_putaddrout2_in = {zll_main_putaddrout7_in[90:85], zll_main_putaddrout7_in[84:0]};
  assign zll_main_putaddrout6_in = {zll_main_putaddrout2_in[90:85], zll_main_putaddrout2_in[84:70]};
  assign zll_main_putaddrout1_in = {zll_main_putaddrout6_in[20:15], zll_main_putaddrout6_in[14:0]};
  assign zll_main_putout12_in = {{zll_main_putaddrout1_in[14], zll_main_putaddrout1_in[20:15], zll_main_putaddrout1_in[7:0]}, zll_main_putaddrout2_in[69:0]};
  ZLL_Main_putOut12  instR1 (zll_main_putout12_in[84:70], zll_main_putout12_in[69:0], zll_main_putout12_out);
  assign res = zll_main_putout12_out;
endmodule

module ZLL_Pure_dispatch7 (input logic [16:0] arg0,
  input logic [69:0] arg1,
  output logic [142:0] res);
  logic [86:0] zll_main_loop220_in;
  logic [86:0] zll_main_putins5_in;
  logic [69:0] zll_main_putins5_out;
  logic [69:0] zll_main_loop226_in;
  logic [142:0] zll_main_loop226_out;
  logic [142:0] zll_main_loop222_in;
  logic [142:0] zll_main_loop222_out;
  assign zll_main_loop220_in = {arg0, arg1};
  assign zll_main_putins5_in = {zll_main_loop220_in[86:70], zll_main_loop220_in[69:0]};
  ZLL_Main_putIns5  inst (zll_main_putins5_in[86:70], zll_main_putins5_in[69:0], zll_main_putins5_out);
  assign zll_main_loop226_in = zll_main_putins5_out;
  ZLL_Main_loop226  instR1 (zll_main_loop226_in[69:0], zll_main_loop226_out);
  assign zll_main_loop222_in = zll_main_loop226_out;
  ZLL_Main_loop222  instR2 (zll_main_loop222_in[142:0], zll_main_loop222_out);
  assign res = zll_main_loop222_out;
endmodule

module ZLL_Main_loop135 (input logic [75:0] arg0,
  output logic [69:0] res);
  logic [75:0] zll_main_finishinstr_in;
  logic [75:0] zll_main_putaddrout4_in;
  logic [69:0] zll_main_putaddrout4_out;
  logic [69:0] main_putweout1_in;
  logic [69:0] main_putweout1_out;
  assign zll_main_finishinstr_in = arg0;
  assign zll_main_putaddrout4_in = {zll_main_finishinstr_in[75:70], zll_main_finishinstr_in[69:0]};
  ZLL_Main_putAddrOut4  inst (zll_main_putaddrout4_in[75:70], zll_main_putaddrout4_in[69:0], zll_main_putaddrout4_out);
  assign main_putweout1_in = zll_main_putaddrout4_out;
  Main_putWeOut1  instR1 (main_putweout1_in[69:0], main_putweout1_out);
  assign res = main_putweout1_out;
endmodule

module ZLL_Main_getReg13 (input logic [1:0] arg0,
  input logic [1:0] arg1,
  input logic [69:0] arg2,
  output logic [77:0] res);
  logic [73:0] zll_main_getreg20_in;
  logic [73:0] zll_main_getreg15_in;
  logic [71:0] zll_main_getreg3_in;
  logic [71:0] zll_main_getreg_in;
  logic [69:0] zll_main_getreg8_in;
  logic [139:0] zll_main_getreg4_in;
  logic [139:0] zll_main_getreg14_in;
  logic [69:0] zll_main_r36_in;
  logic [69:0] zll_main_r3_in;
  logic [61:0] zll_main_r37_in;
  logic [53:0] zll_main_r32_in;
  logic [45:0] zll_main_r35_in;
  logic [7:0] zll_main_r35_out;
  logic [71:0] zll_main_getreg22_in;
  logic [69:0] zll_main_getreg11_in;
  logic [139:0] zll_main_getreg7_in;
  logic [139:0] zll_main_getreg21_in;
  logic [69:0] zll_main_r26_in;
  logic [69:0] zll_main_r21_in;
  logic [61:0] zll_main_r24_in;
  logic [53:0] zll_main_r07_in;
  logic [7:0] zll_main_r07_out;
  logic [71:0] zll_main_getreg5_in;
  logic [69:0] zll_main_getreg18_in;
  logic [139:0] zll_main_getreg1_in;
  logic [139:0] zll_main_getreg16_in;
  logic [69:0] zll_main_r1_in;
  logic [69:0] zll_main_r16_in;
  logic [61:0] zll_main_r17_in;
  logic [7:0] zll_main_r17_out;
  logic [71:0] zll_main_getreg12_in;
  logic [69:0] zll_main_getreg9_in;
  logic [139:0] zll_main_getreg10_in;
  logic [139:0] zll_main_getreg6_in;
  logic [69:0] zll_main_r0_in;
  logic [69:0] zll_main_r02_in;
  logic [61:0] zll_main_r17_inR1;
  logic [7:0] zll_main_r17_outR1;
  assign zll_main_getreg20_in = {arg0, arg0, arg2};
  assign zll_main_getreg15_in = {zll_main_getreg20_in[73:72], zll_main_getreg20_in[73:72], zll_main_getreg20_in[69:0]};
  assign zll_main_getreg3_in = {zll_main_getreg15_in[73:72], zll_main_getreg15_in[69:0]};
  assign zll_main_getreg_in = {zll_main_getreg3_in[69:0], zll_main_getreg3_in[71:70]};
  assign zll_main_getreg8_in = zll_main_getreg_in[71:2];
  assign zll_main_getreg4_in = {zll_main_getreg8_in[69:0], zll_main_getreg8_in[69:0]};
  assign zll_main_getreg14_in = zll_main_getreg4_in[139:0];
  assign zll_main_r36_in = zll_main_getreg14_in[139:70];
  assign zll_main_r3_in = zll_main_r36_in[69:0];
  assign zll_main_r37_in = {zll_main_r3_in[61:54], zll_main_r3_in[53:46], zll_main_r3_in[45:38], zll_main_r3_in[37:32], zll_main_r3_in[31:15], zll_main_r3_in[14:0]};
  assign zll_main_r32_in = {zll_main_r37_in[53:46], zll_main_r37_in[45:38], zll_main_r37_in[37:32], zll_main_r37_in[31:15], zll_main_r37_in[14:0]};
  assign zll_main_r35_in = {zll_main_r32_in[45:38], zll_main_r32_in[37:32], zll_main_r32_in[31:15], zll_main_r32_in[14:0]};
  ZLL_Main_r35  inst (zll_main_r35_in[45:38], zll_main_r35_in[37:32], zll_main_r35_in[31:15], zll_main_r35_in[14:0], zll_main_r35_out);
  assign zll_main_getreg22_in = {zll_main_getreg15_in[69:0], zll_main_getreg15_in[71:70]};
  assign zll_main_getreg11_in = zll_main_getreg22_in[71:2];
  assign zll_main_getreg7_in = {zll_main_getreg11_in[69:0], zll_main_getreg11_in[69:0]};
  assign zll_main_getreg21_in = zll_main_getreg7_in[139:0];
  assign zll_main_r26_in = zll_main_getreg21_in[139:70];
  assign zll_main_r21_in = zll_main_r26_in[69:0];
  assign zll_main_r24_in = {zll_main_r21_in[61:54], zll_main_r21_in[53:46], zll_main_r21_in[45:38], zll_main_r21_in[37:32], zll_main_r21_in[31:15], zll_main_r21_in[14:0]};
  assign zll_main_r07_in = {zll_main_r24_in[53:46], zll_main_r24_in[45:38], zll_main_r24_in[37:32], zll_main_r24_in[31:15], zll_main_r24_in[14:0]};
  ZLL_Main_r07  instR1 (zll_main_r07_in[53:46], zll_main_r07_in[45:38], zll_main_r07_in[37:32], zll_main_r07_in[31:15], zll_main_r07_in[14:0], zll_main_r07_out);
  assign zll_main_getreg5_in = {zll_main_getreg20_in[69:0], zll_main_getreg20_in[71:70]};
  assign zll_main_getreg18_in = zll_main_getreg5_in[71:2];
  assign zll_main_getreg1_in = {zll_main_getreg18_in[69:0], zll_main_getreg18_in[69:0]};
  assign zll_main_getreg16_in = zll_main_getreg1_in[139:0];
  assign zll_main_r1_in = zll_main_getreg16_in[139:70];
  assign zll_main_r16_in = zll_main_r1_in[69:0];
  assign zll_main_r17_in = {zll_main_r16_in[61:54], zll_main_r16_in[53:46], zll_main_r16_in[45:38], zll_main_r16_in[37:32], zll_main_r16_in[31:15], zll_main_r16_in[14:0]};
  ZLL_Main_r17  instR2 (zll_main_r17_in[61:54], zll_main_r17_in[53:46], zll_main_r17_in[45:38], zll_main_r17_in[37:32], zll_main_r17_in[31:15], zll_main_r17_in[14:0], zll_main_r17_out);
  assign zll_main_getreg12_in = {arg2, arg1};
  assign zll_main_getreg9_in = zll_main_getreg12_in[71:2];
  assign zll_main_getreg10_in = {zll_main_getreg9_in[69:0], zll_main_getreg9_in[69:0]};
  assign zll_main_getreg6_in = zll_main_getreg10_in[139:0];
  assign zll_main_r0_in = zll_main_getreg6_in[139:70];
  assign zll_main_r02_in = zll_main_r0_in[69:0];
  assign zll_main_r17_inR1 = {zll_main_r02_in[69:62], zll_main_r02_in[53:46], zll_main_r02_in[45:38], zll_main_r02_in[37:32], zll_main_r02_in[31:15], zll_main_r02_in[14:0]};
  ZLL_Main_r17  instR3 (zll_main_r17_inR1[61:54], zll_main_r17_inR1[53:46], zll_main_r17_inR1[45:38], zll_main_r17_inR1[37:32], zll_main_r17_inR1[31:15], zll_main_r17_inR1[14:0], zll_main_r17_outR1);
  assign res = (zll_main_getreg12_in[1:0] == 2'h0) ? {zll_main_r17_outR1, zll_main_getreg6_in[69:0]} : ((zll_main_getreg5_in[1:0] == 2'h1) ? {zll_main_r17_out, zll_main_getreg16_in[69:0]} : ((zll_main_getreg22_in[1:0] == 2'h2) ? {zll_main_r07_out, zll_main_getreg21_in[69:0]} : {zll_main_r35_out, zll_main_getreg14_in[69:0]}));
endmodule

module Main_getOut (input logic [69:0] arg0,
  output logic [84:0] res);
  logic [139:0] zll_main_getout2_in;
  logic [139:0] zll_main_getout1_in;
  logic [69:0] zll_main_outputs4_in;
  logic [69:0] zll_main_outputs_in;
  logic [61:0] zll_main_outputs5_in;
  logic [53:0] zll_main_outputs3_in;
  logic [45:0] zll_main_outputs6_in;
  logic [37:0] zll_main_outputs7_in;
  logic [31:0] zll_main_outputs1_in;
  assign zll_main_getout2_in = {arg0, arg0};
  assign zll_main_getout1_in = zll_main_getout2_in[139:0];
  assign zll_main_outputs4_in = zll_main_getout1_in[139:70];
  assign zll_main_outputs_in = zll_main_outputs4_in[69:0];
  assign zll_main_outputs5_in = {zll_main_outputs_in[61:54], zll_main_outputs_in[53:46], zll_main_outputs_in[45:38], zll_main_outputs_in[37:32], zll_main_outputs_in[31:15], zll_main_outputs_in[14:0]};
  assign zll_main_outputs3_in = {zll_main_outputs5_in[53:46], zll_main_outputs5_in[45:38], zll_main_outputs5_in[37:32], zll_main_outputs5_in[31:15], zll_main_outputs5_in[14:0]};
  assign zll_main_outputs6_in = {zll_main_outputs3_in[45:38], zll_main_outputs3_in[37:32], zll_main_outputs3_in[31:15], zll_main_outputs3_in[14:0]};
  assign zll_main_outputs7_in = {zll_main_outputs6_in[37:32], zll_main_outputs6_in[31:15], zll_main_outputs6_in[14:0]};
  assign zll_main_outputs1_in = {zll_main_outputs7_in[31:15], zll_main_outputs7_in[14:0]};
  assign res = {zll_main_outputs1_in[14:0], zll_main_getout1_in[69:0]};
endmodule

module Main_putWeOut1 (input logic [69:0] arg0,
  output logic [69:0] res);
  logic [70:0] zll_main_putweout6_in;
  logic [69:0] zll_main_putweout6_out;
  assign zll_main_putweout6_in = {1'h0, arg0};
  ZLL_Main_putWeOut6  inst (zll_main_putweout6_in[70], zll_main_putweout6_in[69:0], zll_main_putweout6_out);
  assign res = zll_main_putweout6_out;
endmodule

module ZLL_Main_putIns5 (input logic [16:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [156:0] zll_main_putins14_in;
  logic [156:0] zll_main_putins_in;
  logic [86:0] zll_main_putins1_in;
  logic [86:0] zll_main_putins11_in;
  logic [86:0] zll_main_putins4_in;
  logic [86:0] zll_main_putins13_in;
  logic [86:0] zll_main_putins10_in;
  logic [86:0] zll_main_putins9_in;
  assign zll_main_putins14_in = {arg0, arg1, arg1};
  assign zll_main_putins_in = {zll_main_putins14_in[156:140], zll_main_putins14_in[139:0]};
  assign zll_main_putins1_in = {zll_main_putins_in[156:140], zll_main_putins_in[139:70]};
  assign zll_main_putins11_in = {zll_main_putins1_in[86:70], zll_main_putins1_in[69:0]};
  assign zll_main_putins4_in = {zll_main_putins11_in[86:70], zll_main_putins11_in[61:54], zll_main_putins11_in[69:62], zll_main_putins11_in[53:46], zll_main_putins11_in[45:38], zll_main_putins11_in[37:32], zll_main_putins11_in[31:15], zll_main_putins11_in[14:0]};
  assign zll_main_putins13_in = {zll_main_putins4_in[53:46], zll_main_putins4_in[86:70], zll_main_putins4_in[69:62], zll_main_putins4_in[61:54], zll_main_putins4_in[45:38], zll_main_putins4_in[37:32], zll_main_putins4_in[31:15], zll_main_putins4_in[14:0]};
  assign zll_main_putins10_in = {zll_main_putins13_in[45:38], zll_main_putins13_in[86:79], zll_main_putins13_in[78:62], zll_main_putins13_in[61:54], zll_main_putins13_in[53:46], zll_main_putins13_in[37:32], zll_main_putins13_in[31:15], zll_main_putins13_in[14:0]};
  assign zll_main_putins9_in = {zll_main_putins10_in[37:32], zll_main_putins10_in[86:79], zll_main_putins10_in[78:71], zll_main_putins10_in[70:54], zll_main_putins10_in[53:46], zll_main_putins10_in[45:38], zll_main_putins10_in[31:15], zll_main_putins10_in[14:0]};
  assign res = {zll_main_putins9_in[39:32], zll_main_putins9_in[47:40], zll_main_putins9_in[72:65], zll_main_putins9_in[80:73], zll_main_putins9_in[86:81], zll_main_putins9_in[64:48], zll_main_putins9_in[14:0]};
endmodule

module ZLL_Main_putReg15 (input logic [7:0] arg0,
  input logic [1:0] arg1,
  input logic [9:0] arg2,
  input logic [69:0] arg3,
  output logic [69:0] res);
  logic [89:0] zll_main_putreg30_in;
  logic [89:0] zll_main_putreg50_in;
  logic [79:0] zll_main_putreg63_in;
  logic [79:0] zll_main_putreg55_in;
  logic [77:0] zll_main_putreg60_in;
  logic [77:0] zll_main_putreg53_in;
  logic [147:0] zll_main_putreg13_in;
  logic [147:0] zll_main_putreg62_in;
  logic [77:0] zll_main_putreg6_in;
  logic [77:0] zll_main_putreg61_in;
  logic [77:0] zll_main_putreg52_in;
  logic [69:0] zll_main_putreg11_in;
  logic [79:0] zll_main_putreg41_in;
  logic [77:0] zll_main_putreg34_in;
  logic [77:0] zll_main_putreg1_in;
  logic [147:0] zll_main_putreg42_in;
  logic [147:0] zll_main_putreg44_in;
  logic [77:0] zll_main_putreg28_in;
  logic [77:0] zll_main_putreg31_in;
  logic [77:0] zll_main_putreg25_in;
  logic [69:0] zll_main_putreg20_in;
  logic [69:0] zll_main_putreg27_in;
  logic [79:0] zll_main_putreg37_in;
  logic [77:0] zll_main_putreg56_in;
  logic [77:0] zll_main_putreg57_in;
  logic [147:0] zll_main_putreg43_in;
  logic [147:0] zll_main_putreg16_in;
  logic [77:0] zll_main_putreg33_in;
  logic [77:0] zll_main_putreg21_in;
  logic [77:0] zll_main_putreg26_in;
  logic [69:0] zll_main_putreg51_in;
  logic [69:0] zll_main_putreg3_in;
  logic [69:0] zll_main_putreg17_in;
  logic [79:0] zll_main_putreg54_in;
  logic [77:0] zll_main_putreg4_in;
  logic [77:0] zll_main_putreg48_in;
  logic [147:0] zll_main_putreg29_in;
  logic [147:0] zll_main_putreg64_in;
  logic [77:0] zll_main_putreg49_in;
  logic [77:0] zll_main_putreg23_in;
  logic [69:0] zll_main_putreg9_in;
  logic [69:0] zll_main_putreg67_in;
  logic [69:0] zll_main_putreg18_in;
  logic [69:0] zll_main_putreg66_in;
  assign zll_main_putreg30_in = {arg0, arg1, arg1, arg0, arg3};
  assign zll_main_putreg50_in = {zll_main_putreg30_in[89:82], zll_main_putreg30_in[81:80], zll_main_putreg30_in[81:80], zll_main_putreg30_in[89:82], zll_main_putreg30_in[69:0]};
  assign zll_main_putreg63_in = {zll_main_putreg50_in[81:80], zll_main_putreg50_in[89:82], zll_main_putreg50_in[69:0]};
  assign zll_main_putreg55_in = {zll_main_putreg63_in[69:0], zll_main_putreg63_in[79:70]};
  assign zll_main_putreg60_in = {zll_main_putreg55_in[79:10], zll_main_putreg55_in[7:0]};
  assign zll_main_putreg53_in = {zll_main_putreg60_in[7:0], zll_main_putreg60_in[77:8]};
  assign zll_main_putreg13_in = {zll_main_putreg53_in[77:70], zll_main_putreg53_in[69:0], zll_main_putreg53_in[69:0]};
  assign zll_main_putreg62_in = {zll_main_putreg13_in[147:140], zll_main_putreg13_in[139:0]};
  assign zll_main_putreg6_in = {zll_main_putreg62_in[147:140], zll_main_putreg62_in[139:70]};
  assign zll_main_putreg61_in = {zll_main_putreg6_in[77:70], zll_main_putreg6_in[69:0]};
  assign zll_main_putreg52_in = {zll_main_putreg61_in[77:70], zll_main_putreg61_in[61:54], zll_main_putreg61_in[69:62], zll_main_putreg61_in[53:46], zll_main_putreg61_in[45:38], zll_main_putreg61_in[37:32], zll_main_putreg61_in[31:15], zll_main_putreg61_in[14:0]};
  assign zll_main_putreg11_in = {zll_main_putreg52_in[77:70], zll_main_putreg52_in[69:62], zll_main_putreg52_in[61:54], zll_main_putreg52_in[53:46], zll_main_putreg52_in[37:32], zll_main_putreg52_in[31:15], zll_main_putreg52_in[14:0]};
  assign zll_main_putreg41_in = {zll_main_putreg50_in[69:0], zll_main_putreg50_in[79:70]};
  assign zll_main_putreg34_in = {zll_main_putreg41_in[79:10], zll_main_putreg41_in[7:0]};
  assign zll_main_putreg1_in = {zll_main_putreg34_in[7:0], zll_main_putreg34_in[77:8]};
  assign zll_main_putreg42_in = {zll_main_putreg1_in[77:70], zll_main_putreg1_in[69:0], zll_main_putreg1_in[69:0]};
  assign zll_main_putreg44_in = {zll_main_putreg42_in[147:140], zll_main_putreg42_in[139:0]};
  assign zll_main_putreg28_in = {zll_main_putreg44_in[147:140], zll_main_putreg44_in[139:70]};
  assign zll_main_putreg31_in = {zll_main_putreg28_in[77:70], zll_main_putreg28_in[69:0]};
  assign zll_main_putreg25_in = {zll_main_putreg31_in[61:54], zll_main_putreg31_in[77:70], zll_main_putreg31_in[69:62], zll_main_putreg31_in[53:46], zll_main_putreg31_in[45:38], zll_main_putreg31_in[37:32], zll_main_putreg31_in[31:15], zll_main_putreg31_in[14:0]};
  assign zll_main_putreg20_in = {zll_main_putreg25_in[77:70], zll_main_putreg25_in[69:62], zll_main_putreg25_in[61:54], zll_main_putreg25_in[45:38], zll_main_putreg25_in[37:32], zll_main_putreg25_in[31:15], zll_main_putreg25_in[14:0]};
  assign zll_main_putreg27_in = {zll_main_putreg20_in[45:38], zll_main_putreg20_in[69:62], zll_main_putreg20_in[61:54], zll_main_putreg20_in[53:46], zll_main_putreg20_in[37:32], zll_main_putreg20_in[31:15], zll_main_putreg20_in[14:0]};
  assign zll_main_putreg37_in = {zll_main_putreg30_in[69:0], zll_main_putreg30_in[79:70]};
  assign zll_main_putreg56_in = {zll_main_putreg37_in[79:10], zll_main_putreg37_in[7:0]};
  assign zll_main_putreg57_in = {zll_main_putreg56_in[7:0], zll_main_putreg56_in[77:8]};
  assign zll_main_putreg43_in = {zll_main_putreg57_in[77:70], zll_main_putreg57_in[69:0], zll_main_putreg57_in[69:0]};
  assign zll_main_putreg16_in = {zll_main_putreg43_in[147:140], zll_main_putreg43_in[139:0]};
  assign zll_main_putreg33_in = {zll_main_putreg16_in[147:140], zll_main_putreg16_in[139:70]};
  assign zll_main_putreg21_in = {zll_main_putreg33_in[77:70], zll_main_putreg33_in[69:0]};
  assign zll_main_putreg26_in = {zll_main_putreg21_in[69:62], zll_main_putreg21_in[77:70], zll_main_putreg21_in[61:54], zll_main_putreg21_in[53:46], zll_main_putreg21_in[45:38], zll_main_putreg21_in[37:32], zll_main_putreg21_in[31:15], zll_main_putreg21_in[14:0]};
  assign zll_main_putreg51_in = {zll_main_putreg26_in[77:70], zll_main_putreg26_in[69:62], zll_main_putreg26_in[53:46], zll_main_putreg26_in[45:38], zll_main_putreg26_in[37:32], zll_main_putreg26_in[31:15], zll_main_putreg26_in[14:0]};
  assign zll_main_putreg3_in = {zll_main_putreg51_in[69:62], zll_main_putreg51_in[45:38], zll_main_putreg51_in[61:54], zll_main_putreg51_in[53:46], zll_main_putreg51_in[37:32], zll_main_putreg51_in[31:15], zll_main_putreg51_in[14:0]};
  assign zll_main_putreg17_in = {zll_main_putreg3_in[37:32], zll_main_putreg3_in[69:62], zll_main_putreg3_in[61:54], zll_main_putreg3_in[53:46], zll_main_putreg3_in[45:38], zll_main_putreg3_in[31:15], zll_main_putreg3_in[14:0]};
  assign zll_main_putreg54_in = {arg3, arg2};
  assign zll_main_putreg4_in = {zll_main_putreg54_in[79:10], zll_main_putreg54_in[7:0]};
  assign zll_main_putreg48_in = {zll_main_putreg4_in[7:0], zll_main_putreg4_in[77:8]};
  assign zll_main_putreg29_in = {zll_main_putreg48_in[77:70], zll_main_putreg48_in[69:0], zll_main_putreg48_in[69:0]};
  assign zll_main_putreg64_in = {zll_main_putreg29_in[147:140], zll_main_putreg29_in[139:0]};
  assign zll_main_putreg49_in = {zll_main_putreg64_in[147:140], zll_main_putreg64_in[139:70]};
  assign zll_main_putreg23_in = {zll_main_putreg49_in[77:70], zll_main_putreg49_in[69:0]};
  assign zll_main_putreg9_in = {zll_main_putreg23_in[77:70], zll_main_putreg23_in[61:54], zll_main_putreg23_in[53:46], zll_main_putreg23_in[45:38], zll_main_putreg23_in[37:32], zll_main_putreg23_in[31:15], zll_main_putreg23_in[14:0]};
  assign zll_main_putreg67_in = {zll_main_putreg9_in[69:62], zll_main_putreg9_in[53:46], zll_main_putreg9_in[61:54], zll_main_putreg9_in[45:38], zll_main_putreg9_in[37:32], zll_main_putreg9_in[31:15], zll_main_putreg9_in[14:0]};
  assign zll_main_putreg18_in = {zll_main_putreg67_in[69:62], zll_main_putreg67_in[45:38], zll_main_putreg67_in[61:54], zll_main_putreg67_in[53:46], zll_main_putreg67_in[37:32], zll_main_putreg67_in[31:15], zll_main_putreg67_in[14:0]};
  assign zll_main_putreg66_in = {zll_main_putreg18_in[37:32], zll_main_putreg18_in[69:62], zll_main_putreg18_in[61:54], zll_main_putreg18_in[53:46], zll_main_putreg18_in[45:38], zll_main_putreg18_in[31:15], zll_main_putreg18_in[14:0]};
  assign res = (zll_main_putreg54_in[9:8] == 2'h0) ? {zll_main_putreg66_in[63:56], zll_main_putreg66_in[39:32], zll_main_putreg66_in[47:40], zll_main_putreg66_in[55:48], zll_main_putreg66_in[69:64], zll_main_putreg66_in[31:15], zll_main_putreg66_in[14:0]} : ((zll_main_putreg37_in[9:8] == 2'h1) ? {zll_main_putreg17_in[63:56], zll_main_putreg17_in[47:40], zll_main_putreg17_in[39:32], zll_main_putreg17_in[55:48], zll_main_putreg17_in[69:64], zll_main_putreg17_in[31:15], zll_main_putreg17_in[14:0]} : ((zll_main_putreg41_in[9:8] == 2'h2) ? {zll_main_putreg27_in[45:38], zll_main_putreg27_in[61:54], zll_main_putreg27_in[53:46], zll_main_putreg27_in[69:62], zll_main_putreg27_in[37:32], zll_main_putreg27_in[31:15], zll_main_putreg27_in[14:0]} : {zll_main_putreg11_in[53:46], zll_main_putreg11_in[61:54], zll_main_putreg11_in[45:38], zll_main_putreg11_in[69:62], zll_main_putreg11_in[37:32], zll_main_putreg11_in[31:15], zll_main_putreg11_in[14:0]}));
endmodule

module Main_incrPC (input logic [69:0] arg0,
  output logic [69:0] res);
  logic [69:0] main_getpc_in;
  logic [75:0] main_getpc_out;
  logic [75:0] zll_main_incrpc1_in;
  logic [75:0] zll_main_incrpc_in;
  logic [11:0] binop_in;
  logic [75:0] zll_main_putpc12_in;
  logic [69:0] zll_main_putpc12_out;
  assign main_getpc_in = arg0;
  Main_getPC  inst (main_getpc_in[69:0], main_getpc_out);
  assign zll_main_incrpc1_in = main_getpc_out;
  assign zll_main_incrpc_in = zll_main_incrpc1_in[75:0];
  assign binop_in = {zll_main_incrpc_in[75:70], 6'h1};
  assign zll_main_putpc12_in = {binop_in[11:6] + binop_in[5:0], zll_main_incrpc_in[69:0]};
  ZLL_Main_putPC12  instR1 (zll_main_putpc12_in[75:70], zll_main_putpc12_in[69:0], zll_main_putpc12_out);
  assign res = zll_main_putpc12_out;
endmodule

module Main_getPC (input logic [69:0] arg0,
  output logic [75:0] res);
  logic [139:0] zll_main_getpc2_in;
  logic [139:0] zll_main_getpc1_in;
  logic [69:0] zll_main_pc_in;
  logic [69:0] zll_main_pc5_in;
  logic [61:0] zll_main_pc6_in;
  logic [53:0] zll_main_pc1_in;
  logic [45:0] zll_main_pc2_in;
  logic [37:0] zll_main_pc4_in;
  logic [20:0] zll_main_pc7_in;
  assign zll_main_getpc2_in = {arg0, arg0};
  assign zll_main_getpc1_in = zll_main_getpc2_in[139:0];
  assign zll_main_pc_in = zll_main_getpc1_in[139:70];
  assign zll_main_pc5_in = zll_main_pc_in[69:0];
  assign zll_main_pc6_in = {zll_main_pc5_in[61:54], zll_main_pc5_in[53:46], zll_main_pc5_in[45:38], zll_main_pc5_in[37:32], zll_main_pc5_in[31:15], zll_main_pc5_in[14:0]};
  assign zll_main_pc1_in = {zll_main_pc6_in[53:46], zll_main_pc6_in[45:38], zll_main_pc6_in[37:32], zll_main_pc6_in[31:15], zll_main_pc6_in[14:0]};
  assign zll_main_pc2_in = {zll_main_pc1_in[45:38], zll_main_pc1_in[37:32], zll_main_pc1_in[31:15], zll_main_pc1_in[14:0]};
  assign zll_main_pc4_in = {zll_main_pc2_in[37:32], zll_main_pc2_in[31:15], zll_main_pc2_in[14:0]};
  assign zll_main_pc7_in = {zll_main_pc4_in[37:32], zll_main_pc4_in[14:0]};
  assign res = {zll_main_pc7_in[20:15], zll_main_getpc1_in[69:0]};
endmodule