module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [99:0] __in0,
  output logic [99:0] __out0,
  output logic [99:0] __out1,
  output logic [99:0] __out2,
  output logic [99:0] __out3);
  logic [99:0] main_dev1_in;
  logic [106:0] zll_main_dev20_in;
  logic [0:0] zll_main_dev20_out;
  logic [106:0] zll_main_dev20_inR1;
  logic [0:0] zll_main_dev20_outR1;
  logic [106:0] zll_main_dev20_inR2;
  logic [0:0] zll_main_dev20_outR2;
  logic [106:0] zll_main_dev20_inR3;
  logic [0:0] zll_main_dev20_outR3;
  logic [106:0] zll_main_dev20_inR4;
  logic [0:0] zll_main_dev20_outR4;
  logic [106:0] zll_main_dev20_inR5;
  logic [0:0] zll_main_dev20_outR5;
  logic [106:0] zll_main_dev20_inR6;
  logic [0:0] zll_main_dev20_outR6;
  logic [106:0] zll_main_dev20_inR7;
  logic [0:0] zll_main_dev20_outR7;
  logic [106:0] zll_main_dev20_inR8;
  logic [0:0] zll_main_dev20_outR8;
  logic [106:0] zll_main_dev20_inR9;
  logic [0:0] zll_main_dev20_outR9;
  logic [106:0] zll_main_dev20_inR10;
  logic [0:0] zll_main_dev20_outR10;
  logic [106:0] zll_main_dev20_inR11;
  logic [0:0] zll_main_dev20_outR11;
  logic [106:0] zll_main_dev20_inR12;
  logic [0:0] zll_main_dev20_outR12;
  logic [106:0] zll_main_dev20_inR13;
  logic [0:0] zll_main_dev20_outR13;
  logic [106:0] zll_main_dev20_inR14;
  logic [0:0] zll_main_dev20_outR14;
  logic [106:0] zll_main_dev20_inR15;
  logic [0:0] zll_main_dev20_outR15;
  logic [106:0] zll_main_dev20_inR16;
  logic [0:0] zll_main_dev20_outR16;
  logic [106:0] zll_main_dev20_inR17;
  logic [0:0] zll_main_dev20_outR17;
  logic [106:0] zll_main_dev20_inR18;
  logic [0:0] zll_main_dev20_outR18;
  logic [106:0] zll_main_dev20_inR19;
  logic [0:0] zll_main_dev20_outR19;
  logic [106:0] zll_main_dev20_inR20;
  logic [0:0] zll_main_dev20_outR20;
  logic [106:0] zll_main_dev20_inR21;
  logic [0:0] zll_main_dev20_outR21;
  logic [106:0] zll_main_dev20_inR22;
  logic [0:0] zll_main_dev20_outR22;
  logic [106:0] zll_main_dev20_inR23;
  logic [0:0] zll_main_dev20_outR23;
  logic [106:0] zll_main_dev20_inR24;
  logic [0:0] zll_main_dev20_outR24;
  logic [106:0] zll_main_dev20_inR25;
  logic [0:0] zll_main_dev20_outR25;
  logic [106:0] zll_main_dev20_inR26;
  logic [0:0] zll_main_dev20_outR26;
  logic [106:0] zll_main_dev20_inR27;
  logic [0:0] zll_main_dev20_outR27;
  logic [106:0] zll_main_dev20_inR28;
  logic [0:0] zll_main_dev20_outR28;
  logic [106:0] zll_main_dev20_inR29;
  logic [0:0] zll_main_dev20_outR29;
  logic [106:0] zll_main_dev20_inR30;
  logic [0:0] zll_main_dev20_outR30;
  logic [106:0] zll_main_dev20_inR31;
  logic [0:0] zll_main_dev20_outR31;
  logic [106:0] zll_main_dev20_inR32;
  logic [0:0] zll_main_dev20_outR32;
  logic [106:0] zll_main_dev20_inR33;
  logic [0:0] zll_main_dev20_outR33;
  logic [106:0] zll_main_dev20_inR34;
  logic [0:0] zll_main_dev20_outR34;
  logic [106:0] zll_main_dev20_inR35;
  logic [0:0] zll_main_dev20_outR35;
  logic [106:0] zll_main_dev20_inR36;
  logic [0:0] zll_main_dev20_outR36;
  logic [106:0] zll_main_dev20_inR37;
  logic [0:0] zll_main_dev20_outR37;
  logic [106:0] zll_main_dev20_inR38;
  logic [0:0] zll_main_dev20_outR38;
  logic [106:0] zll_main_dev20_inR39;
  logic [0:0] zll_main_dev20_outR39;
  logic [106:0] zll_main_dev20_inR40;
  logic [0:0] zll_main_dev20_outR40;
  logic [106:0] zll_main_dev20_inR41;
  logic [0:0] zll_main_dev20_outR41;
  logic [106:0] zll_main_dev20_inR42;
  logic [0:0] zll_main_dev20_outR42;
  logic [106:0] zll_main_dev20_inR43;
  logic [0:0] zll_main_dev20_outR43;
  logic [106:0] zll_main_dev20_inR44;
  logic [0:0] zll_main_dev20_outR44;
  logic [106:0] zll_main_dev20_inR45;
  logic [0:0] zll_main_dev20_outR45;
  logic [106:0] zll_main_dev20_inR46;
  logic [0:0] zll_main_dev20_outR46;
  logic [106:0] zll_main_dev20_inR47;
  logic [0:0] zll_main_dev20_outR47;
  logic [106:0] zll_main_dev20_inR48;
  logic [0:0] zll_main_dev20_outR48;
  logic [106:0] zll_main_dev20_inR49;
  logic [0:0] zll_main_dev20_outR49;
  logic [106:0] zll_main_dev20_inR50;
  logic [0:0] zll_main_dev20_outR50;
  logic [106:0] zll_main_dev20_inR51;
  logic [0:0] zll_main_dev20_outR51;
  logic [106:0] zll_main_dev20_inR52;
  logic [0:0] zll_main_dev20_outR52;
  logic [106:0] zll_main_dev20_inR53;
  logic [0:0] zll_main_dev20_outR53;
  logic [106:0] zll_main_dev20_inR54;
  logic [0:0] zll_main_dev20_outR54;
  logic [106:0] zll_main_dev20_inR55;
  logic [0:0] zll_main_dev20_outR55;
  logic [106:0] zll_main_dev20_inR56;
  logic [0:0] zll_main_dev20_outR56;
  logic [106:0] zll_main_dev20_inR57;
  logic [0:0] zll_main_dev20_outR57;
  logic [106:0] zll_main_dev20_inR58;
  logic [0:0] zll_main_dev20_outR58;
  logic [106:0] zll_main_dev20_inR59;
  logic [0:0] zll_main_dev20_outR59;
  logic [106:0] zll_main_dev20_inR60;
  logic [0:0] zll_main_dev20_outR60;
  logic [106:0] zll_main_dev20_inR61;
  logic [0:0] zll_main_dev20_outR61;
  logic [106:0] zll_main_dev20_inR62;
  logic [0:0] zll_main_dev20_outR62;
  logic [106:0] zll_main_dev20_inR63;
  logic [0:0] zll_main_dev20_outR63;
  logic [106:0] zll_main_dev20_inR64;
  logic [0:0] zll_main_dev20_outR64;
  logic [106:0] zll_main_dev20_inR65;
  logic [0:0] zll_main_dev20_outR65;
  logic [106:0] zll_main_dev20_inR66;
  logic [0:0] zll_main_dev20_outR66;
  logic [106:0] zll_main_dev20_inR67;
  logic [0:0] zll_main_dev20_outR67;
  logic [106:0] zll_main_dev20_inR68;
  logic [0:0] zll_main_dev20_outR68;
  logic [106:0] zll_main_dev20_inR69;
  logic [0:0] zll_main_dev20_outR69;
  logic [106:0] zll_main_dev20_inR70;
  logic [0:0] zll_main_dev20_outR70;
  logic [106:0] zll_main_dev20_inR71;
  logic [0:0] zll_main_dev20_outR71;
  logic [106:0] zll_main_dev20_inR72;
  logic [0:0] zll_main_dev20_outR72;
  logic [106:0] zll_main_dev20_inR73;
  logic [0:0] zll_main_dev20_outR73;
  logic [106:0] zll_main_dev20_inR74;
  logic [0:0] zll_main_dev20_outR74;
  logic [106:0] zll_main_dev20_inR75;
  logic [0:0] zll_main_dev20_outR75;
  logic [106:0] zll_main_dev20_inR76;
  logic [0:0] zll_main_dev20_outR76;
  logic [106:0] zll_main_dev20_inR77;
  logic [0:0] zll_main_dev20_outR77;
  logic [106:0] zll_main_dev20_inR78;
  logic [0:0] zll_main_dev20_outR78;
  logic [106:0] zll_main_dev20_inR79;
  logic [0:0] zll_main_dev20_outR79;
  logic [106:0] zll_main_dev20_inR80;
  logic [0:0] zll_main_dev20_outR80;
  logic [106:0] zll_main_dev20_inR81;
  logic [0:0] zll_main_dev20_outR81;
  logic [106:0] zll_main_dev20_inR82;
  logic [0:0] zll_main_dev20_outR82;
  logic [106:0] zll_main_dev20_inR83;
  logic [0:0] zll_main_dev20_outR83;
  logic [106:0] zll_main_dev20_inR84;
  logic [0:0] zll_main_dev20_outR84;
  logic [106:0] zll_main_dev20_inR85;
  logic [0:0] zll_main_dev20_outR85;
  logic [106:0] zll_main_dev20_inR86;
  logic [0:0] zll_main_dev20_outR86;
  logic [106:0] zll_main_dev20_inR87;
  logic [0:0] zll_main_dev20_outR87;
  logic [106:0] zll_main_dev20_inR88;
  logic [0:0] zll_main_dev20_outR88;
  logic [106:0] zll_main_dev20_inR89;
  logic [0:0] zll_main_dev20_outR89;
  logic [106:0] zll_main_dev20_inR90;
  logic [0:0] zll_main_dev20_outR90;
  logic [106:0] zll_main_dev20_inR91;
  logic [0:0] zll_main_dev20_outR91;
  logic [106:0] zll_main_dev20_inR92;
  logic [0:0] zll_main_dev20_outR92;
  logic [106:0] zll_main_dev20_inR93;
  logic [0:0] zll_main_dev20_outR93;
  logic [106:0] zll_main_dev20_inR94;
  logic [0:0] zll_main_dev20_outR94;
  logic [106:0] zll_main_dev20_inR95;
  logic [0:0] zll_main_dev20_outR95;
  logic [106:0] zll_main_dev20_inR96;
  logic [0:0] zll_main_dev20_outR96;
  logic [106:0] zll_main_dev20_inR97;
  logic [0:0] zll_main_dev20_outR97;
  logic [106:0] zll_main_dev20_inR98;
  logic [0:0] zll_main_dev20_outR98;
  logic [106:0] zll_main_dev20_inR99;
  logic [0:0] zll_main_dev20_outR99;
  logic [106:0] zll_main_dev12_in;
  logic [0:0] zll_main_dev12_out;
  logic [106:0] zll_main_dev12_inR1;
  logic [0:0] zll_main_dev12_outR1;
  logic [106:0] zll_main_dev12_inR2;
  logic [0:0] zll_main_dev12_outR2;
  logic [106:0] zll_main_dev12_inR3;
  logic [0:0] zll_main_dev12_outR3;
  logic [106:0] zll_main_dev12_inR4;
  logic [0:0] zll_main_dev12_outR4;
  logic [106:0] zll_main_dev12_inR5;
  logic [0:0] zll_main_dev12_outR5;
  logic [106:0] zll_main_dev12_inR6;
  logic [0:0] zll_main_dev12_outR6;
  logic [106:0] zll_main_dev12_inR7;
  logic [0:0] zll_main_dev12_outR7;
  logic [106:0] zll_main_dev12_inR8;
  logic [0:0] zll_main_dev12_outR8;
  logic [106:0] zll_main_dev12_inR9;
  logic [0:0] zll_main_dev12_outR9;
  logic [106:0] zll_main_dev12_inR10;
  logic [0:0] zll_main_dev12_outR10;
  logic [106:0] zll_main_dev12_inR11;
  logic [0:0] zll_main_dev12_outR11;
  logic [106:0] zll_main_dev12_inR12;
  logic [0:0] zll_main_dev12_outR12;
  logic [106:0] zll_main_dev12_inR13;
  logic [0:0] zll_main_dev12_outR13;
  logic [106:0] zll_main_dev12_inR14;
  logic [0:0] zll_main_dev12_outR14;
  logic [106:0] zll_main_dev12_inR15;
  logic [0:0] zll_main_dev12_outR15;
  logic [106:0] zll_main_dev12_inR16;
  logic [0:0] zll_main_dev12_outR16;
  logic [106:0] zll_main_dev12_inR17;
  logic [0:0] zll_main_dev12_outR17;
  logic [106:0] zll_main_dev12_inR18;
  logic [0:0] zll_main_dev12_outR18;
  logic [106:0] zll_main_dev12_inR19;
  logic [0:0] zll_main_dev12_outR19;
  logic [106:0] zll_main_dev12_inR20;
  logic [0:0] zll_main_dev12_outR20;
  logic [106:0] zll_main_dev12_inR21;
  logic [0:0] zll_main_dev12_outR21;
  logic [106:0] zll_main_dev12_inR22;
  logic [0:0] zll_main_dev12_outR22;
  logic [106:0] zll_main_dev12_inR23;
  logic [0:0] zll_main_dev12_outR23;
  logic [106:0] zll_main_dev12_inR24;
  logic [0:0] zll_main_dev12_outR24;
  logic [106:0] zll_main_dev12_inR25;
  logic [0:0] zll_main_dev12_outR25;
  logic [106:0] zll_main_dev12_inR26;
  logic [0:0] zll_main_dev12_outR26;
  logic [106:0] zll_main_dev12_inR27;
  logic [0:0] zll_main_dev12_outR27;
  logic [106:0] zll_main_dev12_inR28;
  logic [0:0] zll_main_dev12_outR28;
  logic [106:0] zll_main_dev12_inR29;
  logic [0:0] zll_main_dev12_outR29;
  logic [106:0] zll_main_dev12_inR30;
  logic [0:0] zll_main_dev12_outR30;
  logic [106:0] zll_main_dev12_inR31;
  logic [0:0] zll_main_dev12_outR31;
  logic [106:0] zll_main_dev12_inR32;
  logic [0:0] zll_main_dev12_outR32;
  logic [106:0] zll_main_dev12_inR33;
  logic [0:0] zll_main_dev12_outR33;
  logic [106:0] zll_main_dev12_inR34;
  logic [0:0] zll_main_dev12_outR34;
  logic [106:0] zll_main_dev12_inR35;
  logic [0:0] zll_main_dev12_outR35;
  logic [106:0] zll_main_dev12_inR36;
  logic [0:0] zll_main_dev12_outR36;
  logic [106:0] zll_main_dev12_inR37;
  logic [0:0] zll_main_dev12_outR37;
  logic [106:0] zll_main_dev12_inR38;
  logic [0:0] zll_main_dev12_outR38;
  logic [106:0] zll_main_dev12_inR39;
  logic [0:0] zll_main_dev12_outR39;
  logic [106:0] zll_main_dev12_inR40;
  logic [0:0] zll_main_dev12_outR40;
  logic [106:0] zll_main_dev12_inR41;
  logic [0:0] zll_main_dev12_outR41;
  logic [106:0] zll_main_dev12_inR42;
  logic [0:0] zll_main_dev12_outR42;
  logic [106:0] zll_main_dev12_inR43;
  logic [0:0] zll_main_dev12_outR43;
  logic [106:0] zll_main_dev12_inR44;
  logic [0:0] zll_main_dev12_outR44;
  logic [106:0] zll_main_dev12_inR45;
  logic [0:0] zll_main_dev12_outR45;
  logic [106:0] zll_main_dev12_inR46;
  logic [0:0] zll_main_dev12_outR46;
  logic [106:0] zll_main_dev12_inR47;
  logic [0:0] zll_main_dev12_outR47;
  logic [106:0] zll_main_dev12_inR48;
  logic [0:0] zll_main_dev12_outR48;
  logic [106:0] zll_main_dev12_inR49;
  logic [0:0] zll_main_dev12_outR49;
  logic [106:0] zll_main_dev12_inR50;
  logic [0:0] zll_main_dev12_outR50;
  logic [106:0] zll_main_dev12_inR51;
  logic [0:0] zll_main_dev12_outR51;
  logic [106:0] zll_main_dev12_inR52;
  logic [0:0] zll_main_dev12_outR52;
  logic [106:0] zll_main_dev12_inR53;
  logic [0:0] zll_main_dev12_outR53;
  logic [106:0] zll_main_dev12_inR54;
  logic [0:0] zll_main_dev12_outR54;
  logic [106:0] zll_main_dev12_inR55;
  logic [0:0] zll_main_dev12_outR55;
  logic [106:0] zll_main_dev12_inR56;
  logic [0:0] zll_main_dev12_outR56;
  logic [106:0] zll_main_dev12_inR57;
  logic [0:0] zll_main_dev12_outR57;
  logic [106:0] zll_main_dev12_inR58;
  logic [0:0] zll_main_dev12_outR58;
  logic [106:0] zll_main_dev12_inR59;
  logic [0:0] zll_main_dev12_outR59;
  logic [106:0] zll_main_dev12_inR60;
  logic [0:0] zll_main_dev12_outR60;
  logic [106:0] zll_main_dev12_inR61;
  logic [0:0] zll_main_dev12_outR61;
  logic [106:0] zll_main_dev12_inR62;
  logic [0:0] zll_main_dev12_outR62;
  logic [106:0] zll_main_dev12_inR63;
  logic [0:0] zll_main_dev12_outR63;
  logic [106:0] zll_main_dev12_inR64;
  logic [0:0] zll_main_dev12_outR64;
  logic [106:0] zll_main_dev12_inR65;
  logic [0:0] zll_main_dev12_outR65;
  logic [106:0] zll_main_dev12_inR66;
  logic [0:0] zll_main_dev12_outR66;
  logic [106:0] zll_main_dev12_inR67;
  logic [0:0] zll_main_dev12_outR67;
  logic [106:0] zll_main_dev12_inR68;
  logic [0:0] zll_main_dev12_outR68;
  logic [106:0] zll_main_dev12_inR69;
  logic [0:0] zll_main_dev12_outR69;
  logic [106:0] zll_main_dev12_inR70;
  logic [0:0] zll_main_dev12_outR70;
  logic [106:0] zll_main_dev12_inR71;
  logic [0:0] zll_main_dev12_outR71;
  logic [106:0] zll_main_dev12_inR72;
  logic [0:0] zll_main_dev12_outR72;
  logic [106:0] zll_main_dev12_inR73;
  logic [0:0] zll_main_dev12_outR73;
  logic [106:0] zll_main_dev12_inR74;
  logic [0:0] zll_main_dev12_outR74;
  logic [106:0] zll_main_dev12_inR75;
  logic [0:0] zll_main_dev12_outR75;
  logic [106:0] zll_main_dev12_inR76;
  logic [0:0] zll_main_dev12_outR76;
  logic [106:0] zll_main_dev12_inR77;
  logic [0:0] zll_main_dev12_outR77;
  logic [106:0] zll_main_dev12_inR78;
  logic [0:0] zll_main_dev12_outR78;
  logic [106:0] zll_main_dev12_inR79;
  logic [0:0] zll_main_dev12_outR79;
  logic [106:0] zll_main_dev12_inR80;
  logic [0:0] zll_main_dev12_outR80;
  logic [106:0] zll_main_dev12_inR81;
  logic [0:0] zll_main_dev12_outR81;
  logic [106:0] zll_main_dev12_inR82;
  logic [0:0] zll_main_dev12_outR82;
  logic [106:0] zll_main_dev12_inR83;
  logic [0:0] zll_main_dev12_outR83;
  logic [106:0] zll_main_dev12_inR84;
  logic [0:0] zll_main_dev12_outR84;
  logic [106:0] zll_main_dev12_inR85;
  logic [0:0] zll_main_dev12_outR85;
  logic [106:0] zll_main_dev12_inR86;
  logic [0:0] zll_main_dev12_outR86;
  logic [106:0] zll_main_dev12_inR87;
  logic [0:0] zll_main_dev12_outR87;
  logic [106:0] zll_main_dev12_inR88;
  logic [0:0] zll_main_dev12_outR88;
  logic [106:0] zll_main_dev12_inR89;
  logic [0:0] zll_main_dev12_outR89;
  logic [106:0] zll_main_dev12_inR90;
  logic [0:0] zll_main_dev12_outR90;
  logic [106:0] zll_main_dev12_inR91;
  logic [0:0] zll_main_dev12_outR91;
  logic [106:0] zll_main_dev12_inR92;
  logic [0:0] zll_main_dev12_outR92;
  logic [106:0] zll_main_dev12_inR93;
  logic [0:0] zll_main_dev12_outR93;
  logic [106:0] zll_main_dev12_inR94;
  logic [0:0] zll_main_dev12_outR94;
  logic [106:0] zll_main_dev12_inR95;
  logic [0:0] zll_main_dev12_outR95;
  logic [106:0] zll_main_dev12_inR96;
  logic [0:0] zll_main_dev12_outR96;
  logic [106:0] zll_main_dev12_inR97;
  logic [0:0] zll_main_dev12_outR97;
  logic [106:0] zll_main_dev12_inR98;
  logic [0:0] zll_main_dev12_outR98;
  logic [106:0] zll_main_dev12_inR99;
  logic [0:0] zll_main_dev12_outR99;
  logic [106:0] zll_main_dev15_in;
  logic [0:0] zll_main_dev15_out;
  logic [106:0] zll_main_dev15_inR1;
  logic [0:0] zll_main_dev15_outR1;
  logic [106:0] zll_main_dev15_inR2;
  logic [0:0] zll_main_dev15_outR2;
  logic [106:0] zll_main_dev15_inR3;
  logic [0:0] zll_main_dev15_outR3;
  logic [106:0] zll_main_dev15_inR4;
  logic [0:0] zll_main_dev15_outR4;
  logic [106:0] zll_main_dev15_inR5;
  logic [0:0] zll_main_dev15_outR5;
  logic [106:0] zll_main_dev15_inR6;
  logic [0:0] zll_main_dev15_outR6;
  logic [106:0] zll_main_dev15_inR7;
  logic [0:0] zll_main_dev15_outR7;
  logic [106:0] zll_main_dev15_inR8;
  logic [0:0] zll_main_dev15_outR8;
  logic [106:0] zll_main_dev15_inR9;
  logic [0:0] zll_main_dev15_outR9;
  logic [106:0] zll_main_dev15_inR10;
  logic [0:0] zll_main_dev15_outR10;
  logic [106:0] zll_main_dev15_inR11;
  logic [0:0] zll_main_dev15_outR11;
  logic [106:0] zll_main_dev15_inR12;
  logic [0:0] zll_main_dev15_outR12;
  logic [106:0] zll_main_dev15_inR13;
  logic [0:0] zll_main_dev15_outR13;
  logic [106:0] zll_main_dev15_inR14;
  logic [0:0] zll_main_dev15_outR14;
  logic [106:0] zll_main_dev15_inR15;
  logic [0:0] zll_main_dev15_outR15;
  logic [106:0] zll_main_dev15_inR16;
  logic [0:0] zll_main_dev15_outR16;
  logic [106:0] zll_main_dev15_inR17;
  logic [0:0] zll_main_dev15_outR17;
  logic [106:0] zll_main_dev15_inR18;
  logic [0:0] zll_main_dev15_outR18;
  logic [106:0] zll_main_dev15_inR19;
  logic [0:0] zll_main_dev15_outR19;
  logic [106:0] zll_main_dev15_inR20;
  logic [0:0] zll_main_dev15_outR20;
  logic [106:0] zll_main_dev15_inR21;
  logic [0:0] zll_main_dev15_outR21;
  logic [106:0] zll_main_dev15_inR22;
  logic [0:0] zll_main_dev15_outR22;
  logic [106:0] zll_main_dev15_inR23;
  logic [0:0] zll_main_dev15_outR23;
  logic [106:0] zll_main_dev15_inR24;
  logic [0:0] zll_main_dev15_outR24;
  logic [106:0] zll_main_dev15_inR25;
  logic [0:0] zll_main_dev15_outR25;
  logic [106:0] zll_main_dev15_inR26;
  logic [0:0] zll_main_dev15_outR26;
  logic [106:0] zll_main_dev15_inR27;
  logic [0:0] zll_main_dev15_outR27;
  logic [106:0] zll_main_dev15_inR28;
  logic [0:0] zll_main_dev15_outR28;
  logic [106:0] zll_main_dev15_inR29;
  logic [0:0] zll_main_dev15_outR29;
  logic [106:0] zll_main_dev15_inR30;
  logic [0:0] zll_main_dev15_outR30;
  logic [106:0] zll_main_dev15_inR31;
  logic [0:0] zll_main_dev15_outR31;
  logic [106:0] zll_main_dev15_inR32;
  logic [0:0] zll_main_dev15_outR32;
  logic [106:0] zll_main_dev15_inR33;
  logic [0:0] zll_main_dev15_outR33;
  logic [106:0] zll_main_dev15_inR34;
  logic [0:0] zll_main_dev15_outR34;
  logic [106:0] zll_main_dev15_inR35;
  logic [0:0] zll_main_dev15_outR35;
  logic [106:0] zll_main_dev15_inR36;
  logic [0:0] zll_main_dev15_outR36;
  logic [106:0] zll_main_dev15_inR37;
  logic [0:0] zll_main_dev15_outR37;
  logic [106:0] zll_main_dev15_inR38;
  logic [0:0] zll_main_dev15_outR38;
  logic [106:0] zll_main_dev15_inR39;
  logic [0:0] zll_main_dev15_outR39;
  logic [106:0] zll_main_dev15_inR40;
  logic [0:0] zll_main_dev15_outR40;
  logic [106:0] zll_main_dev15_inR41;
  logic [0:0] zll_main_dev15_outR41;
  logic [106:0] zll_main_dev15_inR42;
  logic [0:0] zll_main_dev15_outR42;
  logic [106:0] zll_main_dev15_inR43;
  logic [0:0] zll_main_dev15_outR43;
  logic [106:0] zll_main_dev15_inR44;
  logic [0:0] zll_main_dev15_outR44;
  logic [106:0] zll_main_dev15_inR45;
  logic [0:0] zll_main_dev15_outR45;
  logic [106:0] zll_main_dev15_inR46;
  logic [0:0] zll_main_dev15_outR46;
  logic [106:0] zll_main_dev15_inR47;
  logic [0:0] zll_main_dev15_outR47;
  logic [106:0] zll_main_dev15_inR48;
  logic [0:0] zll_main_dev15_outR48;
  logic [106:0] zll_main_dev15_inR49;
  logic [0:0] zll_main_dev15_outR49;
  logic [106:0] zll_main_dev15_inR50;
  logic [0:0] zll_main_dev15_outR50;
  logic [106:0] zll_main_dev15_inR51;
  logic [0:0] zll_main_dev15_outR51;
  logic [106:0] zll_main_dev15_inR52;
  logic [0:0] zll_main_dev15_outR52;
  logic [106:0] zll_main_dev15_inR53;
  logic [0:0] zll_main_dev15_outR53;
  logic [106:0] zll_main_dev15_inR54;
  logic [0:0] zll_main_dev15_outR54;
  logic [106:0] zll_main_dev15_inR55;
  logic [0:0] zll_main_dev15_outR55;
  logic [106:0] zll_main_dev15_inR56;
  logic [0:0] zll_main_dev15_outR56;
  logic [106:0] zll_main_dev15_inR57;
  logic [0:0] zll_main_dev15_outR57;
  logic [106:0] zll_main_dev15_inR58;
  logic [0:0] zll_main_dev15_outR58;
  logic [106:0] zll_main_dev15_inR59;
  logic [0:0] zll_main_dev15_outR59;
  logic [106:0] zll_main_dev15_inR60;
  logic [0:0] zll_main_dev15_outR60;
  logic [106:0] zll_main_dev15_inR61;
  logic [0:0] zll_main_dev15_outR61;
  logic [106:0] zll_main_dev15_inR62;
  logic [0:0] zll_main_dev15_outR62;
  logic [106:0] zll_main_dev15_inR63;
  logic [0:0] zll_main_dev15_outR63;
  logic [106:0] zll_main_dev15_inR64;
  logic [0:0] zll_main_dev15_outR64;
  logic [106:0] zll_main_dev15_inR65;
  logic [0:0] zll_main_dev15_outR65;
  logic [106:0] zll_main_dev15_inR66;
  logic [0:0] zll_main_dev15_outR66;
  logic [106:0] zll_main_dev15_inR67;
  logic [0:0] zll_main_dev15_outR67;
  logic [106:0] zll_main_dev15_inR68;
  logic [0:0] zll_main_dev15_outR68;
  logic [106:0] zll_main_dev15_inR69;
  logic [0:0] zll_main_dev15_outR69;
  logic [106:0] zll_main_dev15_inR70;
  logic [0:0] zll_main_dev15_outR70;
  logic [106:0] zll_main_dev15_inR71;
  logic [0:0] zll_main_dev15_outR71;
  logic [106:0] zll_main_dev15_inR72;
  logic [0:0] zll_main_dev15_outR72;
  logic [106:0] zll_main_dev15_inR73;
  logic [0:0] zll_main_dev15_outR73;
  logic [106:0] zll_main_dev15_inR74;
  logic [0:0] zll_main_dev15_outR74;
  logic [106:0] zll_main_dev15_inR75;
  logic [0:0] zll_main_dev15_outR75;
  logic [106:0] zll_main_dev15_inR76;
  logic [0:0] zll_main_dev15_outR76;
  logic [106:0] zll_main_dev15_inR77;
  logic [0:0] zll_main_dev15_outR77;
  logic [106:0] zll_main_dev15_inR78;
  logic [0:0] zll_main_dev15_outR78;
  logic [106:0] zll_main_dev15_inR79;
  logic [0:0] zll_main_dev15_outR79;
  logic [106:0] zll_main_dev15_inR80;
  logic [0:0] zll_main_dev15_outR80;
  logic [106:0] zll_main_dev15_inR81;
  logic [0:0] zll_main_dev15_outR81;
  logic [106:0] zll_main_dev15_inR82;
  logic [0:0] zll_main_dev15_outR82;
  logic [106:0] zll_main_dev15_inR83;
  logic [0:0] zll_main_dev15_outR83;
  logic [106:0] zll_main_dev15_inR84;
  logic [0:0] zll_main_dev15_outR84;
  logic [106:0] zll_main_dev15_inR85;
  logic [0:0] zll_main_dev15_outR85;
  logic [106:0] zll_main_dev15_inR86;
  logic [0:0] zll_main_dev15_outR86;
  logic [106:0] zll_main_dev15_inR87;
  logic [0:0] zll_main_dev15_outR87;
  logic [106:0] zll_main_dev15_inR88;
  logic [0:0] zll_main_dev15_outR88;
  logic [106:0] zll_main_dev15_inR89;
  logic [0:0] zll_main_dev15_outR89;
  logic [106:0] zll_main_dev15_inR90;
  logic [0:0] zll_main_dev15_outR90;
  logic [106:0] zll_main_dev15_inR91;
  logic [0:0] zll_main_dev15_outR91;
  logic [106:0] zll_main_dev15_inR92;
  logic [0:0] zll_main_dev15_outR92;
  logic [106:0] zll_main_dev15_inR93;
  logic [0:0] zll_main_dev15_outR93;
  logic [106:0] zll_main_dev15_inR94;
  logic [0:0] zll_main_dev15_outR94;
  logic [106:0] zll_main_dev15_inR95;
  logic [0:0] zll_main_dev15_outR95;
  logic [106:0] zll_main_dev15_inR96;
  logic [0:0] zll_main_dev15_outR96;
  logic [106:0] zll_main_dev15_inR97;
  logic [0:0] zll_main_dev15_outR97;
  logic [106:0] zll_main_dev15_inR98;
  logic [0:0] zll_main_dev15_outR98;
  logic [106:0] zll_main_dev15_inR99;
  logic [0:0] zll_main_dev15_outR99;
  logic [106:0] zll_main_dev8_in;
  logic [0:0] zll_main_dev8_out;
  logic [106:0] zll_main_dev8_inR1;
  logic [0:0] zll_main_dev8_outR1;
  logic [106:0] zll_main_dev8_inR2;
  logic [0:0] zll_main_dev8_outR2;
  logic [106:0] zll_main_dev8_inR3;
  logic [0:0] zll_main_dev8_outR3;
  logic [106:0] zll_main_dev8_inR4;
  logic [0:0] zll_main_dev8_outR4;
  logic [106:0] zll_main_dev8_inR5;
  logic [0:0] zll_main_dev8_outR5;
  logic [106:0] zll_main_dev8_inR6;
  logic [0:0] zll_main_dev8_outR6;
  logic [106:0] zll_main_dev8_inR7;
  logic [0:0] zll_main_dev8_outR7;
  logic [106:0] zll_main_dev8_inR8;
  logic [0:0] zll_main_dev8_outR8;
  logic [106:0] zll_main_dev8_inR9;
  logic [0:0] zll_main_dev8_outR9;
  logic [106:0] zll_main_dev8_inR10;
  logic [0:0] zll_main_dev8_outR10;
  logic [106:0] zll_main_dev8_inR11;
  logic [0:0] zll_main_dev8_outR11;
  logic [106:0] zll_main_dev8_inR12;
  logic [0:0] zll_main_dev8_outR12;
  logic [106:0] zll_main_dev8_inR13;
  logic [0:0] zll_main_dev8_outR13;
  logic [106:0] zll_main_dev8_inR14;
  logic [0:0] zll_main_dev8_outR14;
  logic [106:0] zll_main_dev8_inR15;
  logic [0:0] zll_main_dev8_outR15;
  logic [106:0] zll_main_dev8_inR16;
  logic [0:0] zll_main_dev8_outR16;
  logic [106:0] zll_main_dev8_inR17;
  logic [0:0] zll_main_dev8_outR17;
  logic [106:0] zll_main_dev8_inR18;
  logic [0:0] zll_main_dev8_outR18;
  logic [106:0] zll_main_dev8_inR19;
  logic [0:0] zll_main_dev8_outR19;
  logic [106:0] zll_main_dev8_inR20;
  logic [0:0] zll_main_dev8_outR20;
  logic [106:0] zll_main_dev8_inR21;
  logic [0:0] zll_main_dev8_outR21;
  logic [106:0] zll_main_dev8_inR22;
  logic [0:0] zll_main_dev8_outR22;
  logic [106:0] zll_main_dev8_inR23;
  logic [0:0] zll_main_dev8_outR23;
  logic [106:0] zll_main_dev8_inR24;
  logic [0:0] zll_main_dev8_outR24;
  logic [106:0] zll_main_dev8_inR25;
  logic [0:0] zll_main_dev8_outR25;
  logic [106:0] zll_main_dev8_inR26;
  logic [0:0] zll_main_dev8_outR26;
  logic [106:0] zll_main_dev8_inR27;
  logic [0:0] zll_main_dev8_outR27;
  logic [106:0] zll_main_dev8_inR28;
  logic [0:0] zll_main_dev8_outR28;
  logic [106:0] zll_main_dev8_inR29;
  logic [0:0] zll_main_dev8_outR29;
  logic [106:0] zll_main_dev8_inR30;
  logic [0:0] zll_main_dev8_outR30;
  logic [106:0] zll_main_dev8_inR31;
  logic [0:0] zll_main_dev8_outR31;
  logic [106:0] zll_main_dev8_inR32;
  logic [0:0] zll_main_dev8_outR32;
  logic [106:0] zll_main_dev8_inR33;
  logic [0:0] zll_main_dev8_outR33;
  logic [106:0] zll_main_dev8_inR34;
  logic [0:0] zll_main_dev8_outR34;
  logic [106:0] zll_main_dev8_inR35;
  logic [0:0] zll_main_dev8_outR35;
  logic [106:0] zll_main_dev8_inR36;
  logic [0:0] zll_main_dev8_outR36;
  logic [106:0] zll_main_dev8_inR37;
  logic [0:0] zll_main_dev8_outR37;
  logic [106:0] zll_main_dev8_inR38;
  logic [0:0] zll_main_dev8_outR38;
  logic [106:0] zll_main_dev8_inR39;
  logic [0:0] zll_main_dev8_outR39;
  logic [106:0] zll_main_dev8_inR40;
  logic [0:0] zll_main_dev8_outR40;
  logic [106:0] zll_main_dev8_inR41;
  logic [0:0] zll_main_dev8_outR41;
  logic [106:0] zll_main_dev8_inR42;
  logic [0:0] zll_main_dev8_outR42;
  logic [106:0] zll_main_dev8_inR43;
  logic [0:0] zll_main_dev8_outR43;
  logic [106:0] zll_main_dev8_inR44;
  logic [0:0] zll_main_dev8_outR44;
  logic [106:0] zll_main_dev8_inR45;
  logic [0:0] zll_main_dev8_outR45;
  logic [106:0] zll_main_dev8_inR46;
  logic [0:0] zll_main_dev8_outR46;
  logic [106:0] zll_main_dev8_inR47;
  logic [0:0] zll_main_dev8_outR47;
  logic [106:0] zll_main_dev8_inR48;
  logic [0:0] zll_main_dev8_outR48;
  logic [106:0] zll_main_dev8_inR49;
  logic [0:0] zll_main_dev8_outR49;
  logic [106:0] zll_main_dev8_inR50;
  logic [0:0] zll_main_dev8_outR50;
  logic [106:0] zll_main_dev8_inR51;
  logic [0:0] zll_main_dev8_outR51;
  logic [106:0] zll_main_dev8_inR52;
  logic [0:0] zll_main_dev8_outR52;
  logic [106:0] zll_main_dev8_inR53;
  logic [0:0] zll_main_dev8_outR53;
  logic [106:0] zll_main_dev8_inR54;
  logic [0:0] zll_main_dev8_outR54;
  logic [106:0] zll_main_dev8_inR55;
  logic [0:0] zll_main_dev8_outR55;
  logic [106:0] zll_main_dev8_inR56;
  logic [0:0] zll_main_dev8_outR56;
  logic [106:0] zll_main_dev8_inR57;
  logic [0:0] zll_main_dev8_outR57;
  logic [106:0] zll_main_dev8_inR58;
  logic [0:0] zll_main_dev8_outR58;
  logic [106:0] zll_main_dev8_inR59;
  logic [0:0] zll_main_dev8_outR59;
  logic [106:0] zll_main_dev8_inR60;
  logic [0:0] zll_main_dev8_outR60;
  logic [106:0] zll_main_dev8_inR61;
  logic [0:0] zll_main_dev8_outR61;
  logic [106:0] zll_main_dev8_inR62;
  logic [0:0] zll_main_dev8_outR62;
  logic [106:0] zll_main_dev8_inR63;
  logic [0:0] zll_main_dev8_outR63;
  logic [106:0] zll_main_dev8_inR64;
  logic [0:0] zll_main_dev8_outR64;
  logic [106:0] zll_main_dev8_inR65;
  logic [0:0] zll_main_dev8_outR65;
  logic [106:0] zll_main_dev8_inR66;
  logic [0:0] zll_main_dev8_outR66;
  logic [106:0] zll_main_dev8_inR67;
  logic [0:0] zll_main_dev8_outR67;
  logic [106:0] zll_main_dev8_inR68;
  logic [0:0] zll_main_dev8_outR68;
  logic [106:0] zll_main_dev8_inR69;
  logic [0:0] zll_main_dev8_outR69;
  logic [106:0] zll_main_dev8_inR70;
  logic [0:0] zll_main_dev8_outR70;
  logic [106:0] zll_main_dev8_inR71;
  logic [0:0] zll_main_dev8_outR71;
  logic [106:0] zll_main_dev8_inR72;
  logic [0:0] zll_main_dev8_outR72;
  logic [106:0] zll_main_dev8_inR73;
  logic [0:0] zll_main_dev8_outR73;
  logic [106:0] zll_main_dev8_inR74;
  logic [0:0] zll_main_dev8_outR74;
  logic [106:0] zll_main_dev8_inR75;
  logic [0:0] zll_main_dev8_outR75;
  logic [106:0] zll_main_dev8_inR76;
  logic [0:0] zll_main_dev8_outR76;
  logic [106:0] zll_main_dev8_inR77;
  logic [0:0] zll_main_dev8_outR77;
  logic [106:0] zll_main_dev8_inR78;
  logic [0:0] zll_main_dev8_outR78;
  logic [106:0] zll_main_dev8_inR79;
  logic [0:0] zll_main_dev8_outR79;
  logic [106:0] zll_main_dev8_inR80;
  logic [0:0] zll_main_dev8_outR80;
  logic [106:0] zll_main_dev8_inR81;
  logic [0:0] zll_main_dev8_outR81;
  logic [106:0] zll_main_dev8_inR82;
  logic [0:0] zll_main_dev8_outR82;
  logic [106:0] zll_main_dev8_inR83;
  logic [0:0] zll_main_dev8_outR83;
  logic [106:0] zll_main_dev8_inR84;
  logic [0:0] zll_main_dev8_outR84;
  logic [106:0] zll_main_dev8_inR85;
  logic [0:0] zll_main_dev8_outR85;
  logic [106:0] zll_main_dev8_inR86;
  logic [0:0] zll_main_dev8_outR86;
  logic [106:0] zll_main_dev8_inR87;
  logic [0:0] zll_main_dev8_outR87;
  logic [106:0] zll_main_dev8_inR88;
  logic [0:0] zll_main_dev8_outR88;
  logic [106:0] zll_main_dev8_inR89;
  logic [0:0] zll_main_dev8_outR89;
  logic [106:0] zll_main_dev8_inR90;
  logic [0:0] zll_main_dev8_outR90;
  logic [106:0] zll_main_dev8_inR91;
  logic [0:0] zll_main_dev8_outR91;
  logic [106:0] zll_main_dev8_inR92;
  logic [0:0] zll_main_dev8_outR92;
  logic [106:0] zll_main_dev8_inR93;
  logic [0:0] zll_main_dev8_outR93;
  logic [106:0] zll_main_dev8_inR94;
  logic [0:0] zll_main_dev8_outR94;
  logic [106:0] zll_main_dev8_inR95;
  logic [0:0] zll_main_dev8_outR95;
  logic [106:0] zll_main_dev8_inR96;
  logic [0:0] zll_main_dev8_outR96;
  logic [106:0] zll_main_dev8_inR97;
  logic [0:0] zll_main_dev8_outR97;
  logic [106:0] zll_main_dev8_inR98;
  logic [0:0] zll_main_dev8_outR98;
  logic [106:0] zll_main_dev8_inR99;
  logic [0:0] zll_main_dev8_outR99;
  logic [0:0] __continue;
  logic [99:0] __resumption_tag;
  logic [99:0] __resumption_tag_next;
  assign main_dev1_in = __resumption_tag;
  assign zll_main_dev20_in = {main_dev1_in[99:0], 7'h0};
  ZLL_Main_dev20  inst (zll_main_dev20_in[106:7], zll_main_dev20_in[6:0], zll_main_dev20_out);
  assign zll_main_dev20_inR1 = {main_dev1_in[99:0], 7'h1};
  ZLL_Main_dev20  instR1 (zll_main_dev20_inR1[106:7], zll_main_dev20_inR1[6:0], zll_main_dev20_outR1);
  assign zll_main_dev20_inR2 = {main_dev1_in[99:0], 7'h2};
  ZLL_Main_dev20  instR2 (zll_main_dev20_inR2[106:7], zll_main_dev20_inR2[6:0], zll_main_dev20_outR2);
  assign zll_main_dev20_inR3 = {main_dev1_in[99:0], 7'h3};
  ZLL_Main_dev20  instR3 (zll_main_dev20_inR3[106:7], zll_main_dev20_inR3[6:0], zll_main_dev20_outR3);
  assign zll_main_dev20_inR4 = {main_dev1_in[99:0], 7'h4};
  ZLL_Main_dev20  instR4 (zll_main_dev20_inR4[106:7], zll_main_dev20_inR4[6:0], zll_main_dev20_outR4);
  assign zll_main_dev20_inR5 = {main_dev1_in[99:0], 7'h5};
  ZLL_Main_dev20  instR5 (zll_main_dev20_inR5[106:7], zll_main_dev20_inR5[6:0], zll_main_dev20_outR5);
  assign zll_main_dev20_inR6 = {main_dev1_in[99:0], 7'h6};
  ZLL_Main_dev20  instR6 (zll_main_dev20_inR6[106:7], zll_main_dev20_inR6[6:0], zll_main_dev20_outR6);
  assign zll_main_dev20_inR7 = {main_dev1_in[99:0], 7'h7};
  ZLL_Main_dev20  instR7 (zll_main_dev20_inR7[106:7], zll_main_dev20_inR7[6:0], zll_main_dev20_outR7);
  assign zll_main_dev20_inR8 = {main_dev1_in[99:0], 7'h8};
  ZLL_Main_dev20  instR8 (zll_main_dev20_inR8[106:7], zll_main_dev20_inR8[6:0], zll_main_dev20_outR8);
  assign zll_main_dev20_inR9 = {main_dev1_in[99:0], 7'h9};
  ZLL_Main_dev20  instR9 (zll_main_dev20_inR9[106:7], zll_main_dev20_inR9[6:0], zll_main_dev20_outR9);
  assign zll_main_dev20_inR10 = {main_dev1_in[99:0], 7'ha};
  ZLL_Main_dev20  instR10 (zll_main_dev20_inR10[106:7], zll_main_dev20_inR10[6:0], zll_main_dev20_outR10);
  assign zll_main_dev20_inR11 = {main_dev1_in[99:0], 7'hb};
  ZLL_Main_dev20  instR11 (zll_main_dev20_inR11[106:7], zll_main_dev20_inR11[6:0], zll_main_dev20_outR11);
  assign zll_main_dev20_inR12 = {main_dev1_in[99:0], 7'hc};
  ZLL_Main_dev20  instR12 (zll_main_dev20_inR12[106:7], zll_main_dev20_inR12[6:0], zll_main_dev20_outR12);
  assign zll_main_dev20_inR13 = {main_dev1_in[99:0], 7'hd};
  ZLL_Main_dev20  instR13 (zll_main_dev20_inR13[106:7], zll_main_dev20_inR13[6:0], zll_main_dev20_outR13);
  assign zll_main_dev20_inR14 = {main_dev1_in[99:0], 7'he};
  ZLL_Main_dev20  instR14 (zll_main_dev20_inR14[106:7], zll_main_dev20_inR14[6:0], zll_main_dev20_outR14);
  assign zll_main_dev20_inR15 = {main_dev1_in[99:0], 7'hf};
  ZLL_Main_dev20  instR15 (zll_main_dev20_inR15[106:7], zll_main_dev20_inR15[6:0], zll_main_dev20_outR15);
  assign zll_main_dev20_inR16 = {main_dev1_in[99:0], 7'h10};
  ZLL_Main_dev20  instR16 (zll_main_dev20_inR16[106:7], zll_main_dev20_inR16[6:0], zll_main_dev20_outR16);
  assign zll_main_dev20_inR17 = {main_dev1_in[99:0], 7'h11};
  ZLL_Main_dev20  instR17 (zll_main_dev20_inR17[106:7], zll_main_dev20_inR17[6:0], zll_main_dev20_outR17);
  assign zll_main_dev20_inR18 = {main_dev1_in[99:0], 7'h12};
  ZLL_Main_dev20  instR18 (zll_main_dev20_inR18[106:7], zll_main_dev20_inR18[6:0], zll_main_dev20_outR18);
  assign zll_main_dev20_inR19 = {main_dev1_in[99:0], 7'h13};
  ZLL_Main_dev20  instR19 (zll_main_dev20_inR19[106:7], zll_main_dev20_inR19[6:0], zll_main_dev20_outR19);
  assign zll_main_dev20_inR20 = {main_dev1_in[99:0], 7'h14};
  ZLL_Main_dev20  instR20 (zll_main_dev20_inR20[106:7], zll_main_dev20_inR20[6:0], zll_main_dev20_outR20);
  assign zll_main_dev20_inR21 = {main_dev1_in[99:0], 7'h15};
  ZLL_Main_dev20  instR21 (zll_main_dev20_inR21[106:7], zll_main_dev20_inR21[6:0], zll_main_dev20_outR21);
  assign zll_main_dev20_inR22 = {main_dev1_in[99:0], 7'h16};
  ZLL_Main_dev20  instR22 (zll_main_dev20_inR22[106:7], zll_main_dev20_inR22[6:0], zll_main_dev20_outR22);
  assign zll_main_dev20_inR23 = {main_dev1_in[99:0], 7'h17};
  ZLL_Main_dev20  instR23 (zll_main_dev20_inR23[106:7], zll_main_dev20_inR23[6:0], zll_main_dev20_outR23);
  assign zll_main_dev20_inR24 = {main_dev1_in[99:0], 7'h18};
  ZLL_Main_dev20  instR24 (zll_main_dev20_inR24[106:7], zll_main_dev20_inR24[6:0], zll_main_dev20_outR24);
  assign zll_main_dev20_inR25 = {main_dev1_in[99:0], 7'h19};
  ZLL_Main_dev20  instR25 (zll_main_dev20_inR25[106:7], zll_main_dev20_inR25[6:0], zll_main_dev20_outR25);
  assign zll_main_dev20_inR26 = {main_dev1_in[99:0], 7'h1a};
  ZLL_Main_dev20  instR26 (zll_main_dev20_inR26[106:7], zll_main_dev20_inR26[6:0], zll_main_dev20_outR26);
  assign zll_main_dev20_inR27 = {main_dev1_in[99:0], 7'h1b};
  ZLL_Main_dev20  instR27 (zll_main_dev20_inR27[106:7], zll_main_dev20_inR27[6:0], zll_main_dev20_outR27);
  assign zll_main_dev20_inR28 = {main_dev1_in[99:0], 7'h1c};
  ZLL_Main_dev20  instR28 (zll_main_dev20_inR28[106:7], zll_main_dev20_inR28[6:0], zll_main_dev20_outR28);
  assign zll_main_dev20_inR29 = {main_dev1_in[99:0], 7'h1d};
  ZLL_Main_dev20  instR29 (zll_main_dev20_inR29[106:7], zll_main_dev20_inR29[6:0], zll_main_dev20_outR29);
  assign zll_main_dev20_inR30 = {main_dev1_in[99:0], 7'h1e};
  ZLL_Main_dev20  instR30 (zll_main_dev20_inR30[106:7], zll_main_dev20_inR30[6:0], zll_main_dev20_outR30);
  assign zll_main_dev20_inR31 = {main_dev1_in[99:0], 7'h1f};
  ZLL_Main_dev20  instR31 (zll_main_dev20_inR31[106:7], zll_main_dev20_inR31[6:0], zll_main_dev20_outR31);
  assign zll_main_dev20_inR32 = {main_dev1_in[99:0], 7'h20};
  ZLL_Main_dev20  instR32 (zll_main_dev20_inR32[106:7], zll_main_dev20_inR32[6:0], zll_main_dev20_outR32);
  assign zll_main_dev20_inR33 = {main_dev1_in[99:0], 7'h21};
  ZLL_Main_dev20  instR33 (zll_main_dev20_inR33[106:7], zll_main_dev20_inR33[6:0], zll_main_dev20_outR33);
  assign zll_main_dev20_inR34 = {main_dev1_in[99:0], 7'h22};
  ZLL_Main_dev20  instR34 (zll_main_dev20_inR34[106:7], zll_main_dev20_inR34[6:0], zll_main_dev20_outR34);
  assign zll_main_dev20_inR35 = {main_dev1_in[99:0], 7'h23};
  ZLL_Main_dev20  instR35 (zll_main_dev20_inR35[106:7], zll_main_dev20_inR35[6:0], zll_main_dev20_outR35);
  assign zll_main_dev20_inR36 = {main_dev1_in[99:0], 7'h24};
  ZLL_Main_dev20  instR36 (zll_main_dev20_inR36[106:7], zll_main_dev20_inR36[6:0], zll_main_dev20_outR36);
  assign zll_main_dev20_inR37 = {main_dev1_in[99:0], 7'h25};
  ZLL_Main_dev20  instR37 (zll_main_dev20_inR37[106:7], zll_main_dev20_inR37[6:0], zll_main_dev20_outR37);
  assign zll_main_dev20_inR38 = {main_dev1_in[99:0], 7'h26};
  ZLL_Main_dev20  instR38 (zll_main_dev20_inR38[106:7], zll_main_dev20_inR38[6:0], zll_main_dev20_outR38);
  assign zll_main_dev20_inR39 = {main_dev1_in[99:0], 7'h27};
  ZLL_Main_dev20  instR39 (zll_main_dev20_inR39[106:7], zll_main_dev20_inR39[6:0], zll_main_dev20_outR39);
  assign zll_main_dev20_inR40 = {main_dev1_in[99:0], 7'h28};
  ZLL_Main_dev20  instR40 (zll_main_dev20_inR40[106:7], zll_main_dev20_inR40[6:0], zll_main_dev20_outR40);
  assign zll_main_dev20_inR41 = {main_dev1_in[99:0], 7'h29};
  ZLL_Main_dev20  instR41 (zll_main_dev20_inR41[106:7], zll_main_dev20_inR41[6:0], zll_main_dev20_outR41);
  assign zll_main_dev20_inR42 = {main_dev1_in[99:0], 7'h2a};
  ZLL_Main_dev20  instR42 (zll_main_dev20_inR42[106:7], zll_main_dev20_inR42[6:0], zll_main_dev20_outR42);
  assign zll_main_dev20_inR43 = {main_dev1_in[99:0], 7'h2b};
  ZLL_Main_dev20  instR43 (zll_main_dev20_inR43[106:7], zll_main_dev20_inR43[6:0], zll_main_dev20_outR43);
  assign zll_main_dev20_inR44 = {main_dev1_in[99:0], 7'h2c};
  ZLL_Main_dev20  instR44 (zll_main_dev20_inR44[106:7], zll_main_dev20_inR44[6:0], zll_main_dev20_outR44);
  assign zll_main_dev20_inR45 = {main_dev1_in[99:0], 7'h2d};
  ZLL_Main_dev20  instR45 (zll_main_dev20_inR45[106:7], zll_main_dev20_inR45[6:0], zll_main_dev20_outR45);
  assign zll_main_dev20_inR46 = {main_dev1_in[99:0], 7'h2e};
  ZLL_Main_dev20  instR46 (zll_main_dev20_inR46[106:7], zll_main_dev20_inR46[6:0], zll_main_dev20_outR46);
  assign zll_main_dev20_inR47 = {main_dev1_in[99:0], 7'h2f};
  ZLL_Main_dev20  instR47 (zll_main_dev20_inR47[106:7], zll_main_dev20_inR47[6:0], zll_main_dev20_outR47);
  assign zll_main_dev20_inR48 = {main_dev1_in[99:0], 7'h30};
  ZLL_Main_dev20  instR48 (zll_main_dev20_inR48[106:7], zll_main_dev20_inR48[6:0], zll_main_dev20_outR48);
  assign zll_main_dev20_inR49 = {main_dev1_in[99:0], 7'h31};
  ZLL_Main_dev20  instR49 (zll_main_dev20_inR49[106:7], zll_main_dev20_inR49[6:0], zll_main_dev20_outR49);
  assign zll_main_dev20_inR50 = {main_dev1_in[99:0], 7'h32};
  ZLL_Main_dev20  instR50 (zll_main_dev20_inR50[106:7], zll_main_dev20_inR50[6:0], zll_main_dev20_outR50);
  assign zll_main_dev20_inR51 = {main_dev1_in[99:0], 7'h33};
  ZLL_Main_dev20  instR51 (zll_main_dev20_inR51[106:7], zll_main_dev20_inR51[6:0], zll_main_dev20_outR51);
  assign zll_main_dev20_inR52 = {main_dev1_in[99:0], 7'h34};
  ZLL_Main_dev20  instR52 (zll_main_dev20_inR52[106:7], zll_main_dev20_inR52[6:0], zll_main_dev20_outR52);
  assign zll_main_dev20_inR53 = {main_dev1_in[99:0], 7'h35};
  ZLL_Main_dev20  instR53 (zll_main_dev20_inR53[106:7], zll_main_dev20_inR53[6:0], zll_main_dev20_outR53);
  assign zll_main_dev20_inR54 = {main_dev1_in[99:0], 7'h36};
  ZLL_Main_dev20  instR54 (zll_main_dev20_inR54[106:7], zll_main_dev20_inR54[6:0], zll_main_dev20_outR54);
  assign zll_main_dev20_inR55 = {main_dev1_in[99:0], 7'h37};
  ZLL_Main_dev20  instR55 (zll_main_dev20_inR55[106:7], zll_main_dev20_inR55[6:0], zll_main_dev20_outR55);
  assign zll_main_dev20_inR56 = {main_dev1_in[99:0], 7'h38};
  ZLL_Main_dev20  instR56 (zll_main_dev20_inR56[106:7], zll_main_dev20_inR56[6:0], zll_main_dev20_outR56);
  assign zll_main_dev20_inR57 = {main_dev1_in[99:0], 7'h39};
  ZLL_Main_dev20  instR57 (zll_main_dev20_inR57[106:7], zll_main_dev20_inR57[6:0], zll_main_dev20_outR57);
  assign zll_main_dev20_inR58 = {main_dev1_in[99:0], 7'h3a};
  ZLL_Main_dev20  instR58 (zll_main_dev20_inR58[106:7], zll_main_dev20_inR58[6:0], zll_main_dev20_outR58);
  assign zll_main_dev20_inR59 = {main_dev1_in[99:0], 7'h3b};
  ZLL_Main_dev20  instR59 (zll_main_dev20_inR59[106:7], zll_main_dev20_inR59[6:0], zll_main_dev20_outR59);
  assign zll_main_dev20_inR60 = {main_dev1_in[99:0], 7'h3c};
  ZLL_Main_dev20  instR60 (zll_main_dev20_inR60[106:7], zll_main_dev20_inR60[6:0], zll_main_dev20_outR60);
  assign zll_main_dev20_inR61 = {main_dev1_in[99:0], 7'h3d};
  ZLL_Main_dev20  instR61 (zll_main_dev20_inR61[106:7], zll_main_dev20_inR61[6:0], zll_main_dev20_outR61);
  assign zll_main_dev20_inR62 = {main_dev1_in[99:0], 7'h3e};
  ZLL_Main_dev20  instR62 (zll_main_dev20_inR62[106:7], zll_main_dev20_inR62[6:0], zll_main_dev20_outR62);
  assign zll_main_dev20_inR63 = {main_dev1_in[99:0], 7'h3f};
  ZLL_Main_dev20  instR63 (zll_main_dev20_inR63[106:7], zll_main_dev20_inR63[6:0], zll_main_dev20_outR63);
  assign zll_main_dev20_inR64 = {main_dev1_in[99:0], 7'h40};
  ZLL_Main_dev20  instR64 (zll_main_dev20_inR64[106:7], zll_main_dev20_inR64[6:0], zll_main_dev20_outR64);
  assign zll_main_dev20_inR65 = {main_dev1_in[99:0], 7'h41};
  ZLL_Main_dev20  instR65 (zll_main_dev20_inR65[106:7], zll_main_dev20_inR65[6:0], zll_main_dev20_outR65);
  assign zll_main_dev20_inR66 = {main_dev1_in[99:0], 7'h42};
  ZLL_Main_dev20  instR66 (zll_main_dev20_inR66[106:7], zll_main_dev20_inR66[6:0], zll_main_dev20_outR66);
  assign zll_main_dev20_inR67 = {main_dev1_in[99:0], 7'h43};
  ZLL_Main_dev20  instR67 (zll_main_dev20_inR67[106:7], zll_main_dev20_inR67[6:0], zll_main_dev20_outR67);
  assign zll_main_dev20_inR68 = {main_dev1_in[99:0], 7'h44};
  ZLL_Main_dev20  instR68 (zll_main_dev20_inR68[106:7], zll_main_dev20_inR68[6:0], zll_main_dev20_outR68);
  assign zll_main_dev20_inR69 = {main_dev1_in[99:0], 7'h45};
  ZLL_Main_dev20  instR69 (zll_main_dev20_inR69[106:7], zll_main_dev20_inR69[6:0], zll_main_dev20_outR69);
  assign zll_main_dev20_inR70 = {main_dev1_in[99:0], 7'h46};
  ZLL_Main_dev20  instR70 (zll_main_dev20_inR70[106:7], zll_main_dev20_inR70[6:0], zll_main_dev20_outR70);
  assign zll_main_dev20_inR71 = {main_dev1_in[99:0], 7'h47};
  ZLL_Main_dev20  instR71 (zll_main_dev20_inR71[106:7], zll_main_dev20_inR71[6:0], zll_main_dev20_outR71);
  assign zll_main_dev20_inR72 = {main_dev1_in[99:0], 7'h48};
  ZLL_Main_dev20  instR72 (zll_main_dev20_inR72[106:7], zll_main_dev20_inR72[6:0], zll_main_dev20_outR72);
  assign zll_main_dev20_inR73 = {main_dev1_in[99:0], 7'h49};
  ZLL_Main_dev20  instR73 (zll_main_dev20_inR73[106:7], zll_main_dev20_inR73[6:0], zll_main_dev20_outR73);
  assign zll_main_dev20_inR74 = {main_dev1_in[99:0], 7'h4a};
  ZLL_Main_dev20  instR74 (zll_main_dev20_inR74[106:7], zll_main_dev20_inR74[6:0], zll_main_dev20_outR74);
  assign zll_main_dev20_inR75 = {main_dev1_in[99:0], 7'h4b};
  ZLL_Main_dev20  instR75 (zll_main_dev20_inR75[106:7], zll_main_dev20_inR75[6:0], zll_main_dev20_outR75);
  assign zll_main_dev20_inR76 = {main_dev1_in[99:0], 7'h4c};
  ZLL_Main_dev20  instR76 (zll_main_dev20_inR76[106:7], zll_main_dev20_inR76[6:0], zll_main_dev20_outR76);
  assign zll_main_dev20_inR77 = {main_dev1_in[99:0], 7'h4d};
  ZLL_Main_dev20  instR77 (zll_main_dev20_inR77[106:7], zll_main_dev20_inR77[6:0], zll_main_dev20_outR77);
  assign zll_main_dev20_inR78 = {main_dev1_in[99:0], 7'h4e};
  ZLL_Main_dev20  instR78 (zll_main_dev20_inR78[106:7], zll_main_dev20_inR78[6:0], zll_main_dev20_outR78);
  assign zll_main_dev20_inR79 = {main_dev1_in[99:0], 7'h4f};
  ZLL_Main_dev20  instR79 (zll_main_dev20_inR79[106:7], zll_main_dev20_inR79[6:0], zll_main_dev20_outR79);
  assign zll_main_dev20_inR80 = {main_dev1_in[99:0], 7'h50};
  ZLL_Main_dev20  instR80 (zll_main_dev20_inR80[106:7], zll_main_dev20_inR80[6:0], zll_main_dev20_outR80);
  assign zll_main_dev20_inR81 = {main_dev1_in[99:0], 7'h51};
  ZLL_Main_dev20  instR81 (zll_main_dev20_inR81[106:7], zll_main_dev20_inR81[6:0], zll_main_dev20_outR81);
  assign zll_main_dev20_inR82 = {main_dev1_in[99:0], 7'h52};
  ZLL_Main_dev20  instR82 (zll_main_dev20_inR82[106:7], zll_main_dev20_inR82[6:0], zll_main_dev20_outR82);
  assign zll_main_dev20_inR83 = {main_dev1_in[99:0], 7'h53};
  ZLL_Main_dev20  instR83 (zll_main_dev20_inR83[106:7], zll_main_dev20_inR83[6:0], zll_main_dev20_outR83);
  assign zll_main_dev20_inR84 = {main_dev1_in[99:0], 7'h54};
  ZLL_Main_dev20  instR84 (zll_main_dev20_inR84[106:7], zll_main_dev20_inR84[6:0], zll_main_dev20_outR84);
  assign zll_main_dev20_inR85 = {main_dev1_in[99:0], 7'h55};
  ZLL_Main_dev20  instR85 (zll_main_dev20_inR85[106:7], zll_main_dev20_inR85[6:0], zll_main_dev20_outR85);
  assign zll_main_dev20_inR86 = {main_dev1_in[99:0], 7'h56};
  ZLL_Main_dev20  instR86 (zll_main_dev20_inR86[106:7], zll_main_dev20_inR86[6:0], zll_main_dev20_outR86);
  assign zll_main_dev20_inR87 = {main_dev1_in[99:0], 7'h57};
  ZLL_Main_dev20  instR87 (zll_main_dev20_inR87[106:7], zll_main_dev20_inR87[6:0], zll_main_dev20_outR87);
  assign zll_main_dev20_inR88 = {main_dev1_in[99:0], 7'h58};
  ZLL_Main_dev20  instR88 (zll_main_dev20_inR88[106:7], zll_main_dev20_inR88[6:0], zll_main_dev20_outR88);
  assign zll_main_dev20_inR89 = {main_dev1_in[99:0], 7'h59};
  ZLL_Main_dev20  instR89 (zll_main_dev20_inR89[106:7], zll_main_dev20_inR89[6:0], zll_main_dev20_outR89);
  assign zll_main_dev20_inR90 = {main_dev1_in[99:0], 7'h5a};
  ZLL_Main_dev20  instR90 (zll_main_dev20_inR90[106:7], zll_main_dev20_inR90[6:0], zll_main_dev20_outR90);
  assign zll_main_dev20_inR91 = {main_dev1_in[99:0], 7'h5b};
  ZLL_Main_dev20  instR91 (zll_main_dev20_inR91[106:7], zll_main_dev20_inR91[6:0], zll_main_dev20_outR91);
  assign zll_main_dev20_inR92 = {main_dev1_in[99:0], 7'h5c};
  ZLL_Main_dev20  instR92 (zll_main_dev20_inR92[106:7], zll_main_dev20_inR92[6:0], zll_main_dev20_outR92);
  assign zll_main_dev20_inR93 = {main_dev1_in[99:0], 7'h5d};
  ZLL_Main_dev20  instR93 (zll_main_dev20_inR93[106:7], zll_main_dev20_inR93[6:0], zll_main_dev20_outR93);
  assign zll_main_dev20_inR94 = {main_dev1_in[99:0], 7'h5e};
  ZLL_Main_dev20  instR94 (zll_main_dev20_inR94[106:7], zll_main_dev20_inR94[6:0], zll_main_dev20_outR94);
  assign zll_main_dev20_inR95 = {main_dev1_in[99:0], 7'h5f};
  ZLL_Main_dev20  instR95 (zll_main_dev20_inR95[106:7], zll_main_dev20_inR95[6:0], zll_main_dev20_outR95);
  assign zll_main_dev20_inR96 = {main_dev1_in[99:0], 7'h60};
  ZLL_Main_dev20  instR96 (zll_main_dev20_inR96[106:7], zll_main_dev20_inR96[6:0], zll_main_dev20_outR96);
  assign zll_main_dev20_inR97 = {main_dev1_in[99:0], 7'h61};
  ZLL_Main_dev20  instR97 (zll_main_dev20_inR97[106:7], zll_main_dev20_inR97[6:0], zll_main_dev20_outR97);
  assign zll_main_dev20_inR98 = {main_dev1_in[99:0], 7'h62};
  ZLL_Main_dev20  instR98 (zll_main_dev20_inR98[106:7], zll_main_dev20_inR98[6:0], zll_main_dev20_outR98);
  assign zll_main_dev20_inR99 = {main_dev1_in[99:0], 7'h63};
  ZLL_Main_dev20  instR99 (zll_main_dev20_inR99[106:7], zll_main_dev20_inR99[6:0], zll_main_dev20_outR99);
  assign zll_main_dev12_in = {main_dev1_in[99:0], 7'h0};
  ZLL_Main_dev12  instR100 (zll_main_dev12_in[106:7], zll_main_dev12_in[6:0], zll_main_dev12_out);
  assign zll_main_dev12_inR1 = {main_dev1_in[99:0], 7'h1};
  ZLL_Main_dev12  instR101 (zll_main_dev12_inR1[106:7], zll_main_dev12_inR1[6:0], zll_main_dev12_outR1);
  assign zll_main_dev12_inR2 = {main_dev1_in[99:0], 7'h2};
  ZLL_Main_dev12  instR102 (zll_main_dev12_inR2[106:7], zll_main_dev12_inR2[6:0], zll_main_dev12_outR2);
  assign zll_main_dev12_inR3 = {main_dev1_in[99:0], 7'h3};
  ZLL_Main_dev12  instR103 (zll_main_dev12_inR3[106:7], zll_main_dev12_inR3[6:0], zll_main_dev12_outR3);
  assign zll_main_dev12_inR4 = {main_dev1_in[99:0], 7'h4};
  ZLL_Main_dev12  instR104 (zll_main_dev12_inR4[106:7], zll_main_dev12_inR4[6:0], zll_main_dev12_outR4);
  assign zll_main_dev12_inR5 = {main_dev1_in[99:0], 7'h5};
  ZLL_Main_dev12  instR105 (zll_main_dev12_inR5[106:7], zll_main_dev12_inR5[6:0], zll_main_dev12_outR5);
  assign zll_main_dev12_inR6 = {main_dev1_in[99:0], 7'h6};
  ZLL_Main_dev12  instR106 (zll_main_dev12_inR6[106:7], zll_main_dev12_inR6[6:0], zll_main_dev12_outR6);
  assign zll_main_dev12_inR7 = {main_dev1_in[99:0], 7'h7};
  ZLL_Main_dev12  instR107 (zll_main_dev12_inR7[106:7], zll_main_dev12_inR7[6:0], zll_main_dev12_outR7);
  assign zll_main_dev12_inR8 = {main_dev1_in[99:0], 7'h8};
  ZLL_Main_dev12  instR108 (zll_main_dev12_inR8[106:7], zll_main_dev12_inR8[6:0], zll_main_dev12_outR8);
  assign zll_main_dev12_inR9 = {main_dev1_in[99:0], 7'h9};
  ZLL_Main_dev12  instR109 (zll_main_dev12_inR9[106:7], zll_main_dev12_inR9[6:0], zll_main_dev12_outR9);
  assign zll_main_dev12_inR10 = {main_dev1_in[99:0], 7'ha};
  ZLL_Main_dev12  instR110 (zll_main_dev12_inR10[106:7], zll_main_dev12_inR10[6:0], zll_main_dev12_outR10);
  assign zll_main_dev12_inR11 = {main_dev1_in[99:0], 7'hb};
  ZLL_Main_dev12  instR111 (zll_main_dev12_inR11[106:7], zll_main_dev12_inR11[6:0], zll_main_dev12_outR11);
  assign zll_main_dev12_inR12 = {main_dev1_in[99:0], 7'hc};
  ZLL_Main_dev12  instR112 (zll_main_dev12_inR12[106:7], zll_main_dev12_inR12[6:0], zll_main_dev12_outR12);
  assign zll_main_dev12_inR13 = {main_dev1_in[99:0], 7'hd};
  ZLL_Main_dev12  instR113 (zll_main_dev12_inR13[106:7], zll_main_dev12_inR13[6:0], zll_main_dev12_outR13);
  assign zll_main_dev12_inR14 = {main_dev1_in[99:0], 7'he};
  ZLL_Main_dev12  instR114 (zll_main_dev12_inR14[106:7], zll_main_dev12_inR14[6:0], zll_main_dev12_outR14);
  assign zll_main_dev12_inR15 = {main_dev1_in[99:0], 7'hf};
  ZLL_Main_dev12  instR115 (zll_main_dev12_inR15[106:7], zll_main_dev12_inR15[6:0], zll_main_dev12_outR15);
  assign zll_main_dev12_inR16 = {main_dev1_in[99:0], 7'h10};
  ZLL_Main_dev12  instR116 (zll_main_dev12_inR16[106:7], zll_main_dev12_inR16[6:0], zll_main_dev12_outR16);
  assign zll_main_dev12_inR17 = {main_dev1_in[99:0], 7'h11};
  ZLL_Main_dev12  instR117 (zll_main_dev12_inR17[106:7], zll_main_dev12_inR17[6:0], zll_main_dev12_outR17);
  assign zll_main_dev12_inR18 = {main_dev1_in[99:0], 7'h12};
  ZLL_Main_dev12  instR118 (zll_main_dev12_inR18[106:7], zll_main_dev12_inR18[6:0], zll_main_dev12_outR18);
  assign zll_main_dev12_inR19 = {main_dev1_in[99:0], 7'h13};
  ZLL_Main_dev12  instR119 (zll_main_dev12_inR19[106:7], zll_main_dev12_inR19[6:0], zll_main_dev12_outR19);
  assign zll_main_dev12_inR20 = {main_dev1_in[99:0], 7'h14};
  ZLL_Main_dev12  instR120 (zll_main_dev12_inR20[106:7], zll_main_dev12_inR20[6:0], zll_main_dev12_outR20);
  assign zll_main_dev12_inR21 = {main_dev1_in[99:0], 7'h15};
  ZLL_Main_dev12  instR121 (zll_main_dev12_inR21[106:7], zll_main_dev12_inR21[6:0], zll_main_dev12_outR21);
  assign zll_main_dev12_inR22 = {main_dev1_in[99:0], 7'h16};
  ZLL_Main_dev12  instR122 (zll_main_dev12_inR22[106:7], zll_main_dev12_inR22[6:0], zll_main_dev12_outR22);
  assign zll_main_dev12_inR23 = {main_dev1_in[99:0], 7'h17};
  ZLL_Main_dev12  instR123 (zll_main_dev12_inR23[106:7], zll_main_dev12_inR23[6:0], zll_main_dev12_outR23);
  assign zll_main_dev12_inR24 = {main_dev1_in[99:0], 7'h18};
  ZLL_Main_dev12  instR124 (zll_main_dev12_inR24[106:7], zll_main_dev12_inR24[6:0], zll_main_dev12_outR24);
  assign zll_main_dev12_inR25 = {main_dev1_in[99:0], 7'h19};
  ZLL_Main_dev12  instR125 (zll_main_dev12_inR25[106:7], zll_main_dev12_inR25[6:0], zll_main_dev12_outR25);
  assign zll_main_dev12_inR26 = {main_dev1_in[99:0], 7'h1a};
  ZLL_Main_dev12  instR126 (zll_main_dev12_inR26[106:7], zll_main_dev12_inR26[6:0], zll_main_dev12_outR26);
  assign zll_main_dev12_inR27 = {main_dev1_in[99:0], 7'h1b};
  ZLL_Main_dev12  instR127 (zll_main_dev12_inR27[106:7], zll_main_dev12_inR27[6:0], zll_main_dev12_outR27);
  assign zll_main_dev12_inR28 = {main_dev1_in[99:0], 7'h1c};
  ZLL_Main_dev12  instR128 (zll_main_dev12_inR28[106:7], zll_main_dev12_inR28[6:0], zll_main_dev12_outR28);
  assign zll_main_dev12_inR29 = {main_dev1_in[99:0], 7'h1d};
  ZLL_Main_dev12  instR129 (zll_main_dev12_inR29[106:7], zll_main_dev12_inR29[6:0], zll_main_dev12_outR29);
  assign zll_main_dev12_inR30 = {main_dev1_in[99:0], 7'h1e};
  ZLL_Main_dev12  instR130 (zll_main_dev12_inR30[106:7], zll_main_dev12_inR30[6:0], zll_main_dev12_outR30);
  assign zll_main_dev12_inR31 = {main_dev1_in[99:0], 7'h1f};
  ZLL_Main_dev12  instR131 (zll_main_dev12_inR31[106:7], zll_main_dev12_inR31[6:0], zll_main_dev12_outR31);
  assign zll_main_dev12_inR32 = {main_dev1_in[99:0], 7'h20};
  ZLL_Main_dev12  instR132 (zll_main_dev12_inR32[106:7], zll_main_dev12_inR32[6:0], zll_main_dev12_outR32);
  assign zll_main_dev12_inR33 = {main_dev1_in[99:0], 7'h21};
  ZLL_Main_dev12  instR133 (zll_main_dev12_inR33[106:7], zll_main_dev12_inR33[6:0], zll_main_dev12_outR33);
  assign zll_main_dev12_inR34 = {main_dev1_in[99:0], 7'h22};
  ZLL_Main_dev12  instR134 (zll_main_dev12_inR34[106:7], zll_main_dev12_inR34[6:0], zll_main_dev12_outR34);
  assign zll_main_dev12_inR35 = {main_dev1_in[99:0], 7'h23};
  ZLL_Main_dev12  instR135 (zll_main_dev12_inR35[106:7], zll_main_dev12_inR35[6:0], zll_main_dev12_outR35);
  assign zll_main_dev12_inR36 = {main_dev1_in[99:0], 7'h24};
  ZLL_Main_dev12  instR136 (zll_main_dev12_inR36[106:7], zll_main_dev12_inR36[6:0], zll_main_dev12_outR36);
  assign zll_main_dev12_inR37 = {main_dev1_in[99:0], 7'h25};
  ZLL_Main_dev12  instR137 (zll_main_dev12_inR37[106:7], zll_main_dev12_inR37[6:0], zll_main_dev12_outR37);
  assign zll_main_dev12_inR38 = {main_dev1_in[99:0], 7'h26};
  ZLL_Main_dev12  instR138 (zll_main_dev12_inR38[106:7], zll_main_dev12_inR38[6:0], zll_main_dev12_outR38);
  assign zll_main_dev12_inR39 = {main_dev1_in[99:0], 7'h27};
  ZLL_Main_dev12  instR139 (zll_main_dev12_inR39[106:7], zll_main_dev12_inR39[6:0], zll_main_dev12_outR39);
  assign zll_main_dev12_inR40 = {main_dev1_in[99:0], 7'h28};
  ZLL_Main_dev12  instR140 (zll_main_dev12_inR40[106:7], zll_main_dev12_inR40[6:0], zll_main_dev12_outR40);
  assign zll_main_dev12_inR41 = {main_dev1_in[99:0], 7'h29};
  ZLL_Main_dev12  instR141 (zll_main_dev12_inR41[106:7], zll_main_dev12_inR41[6:0], zll_main_dev12_outR41);
  assign zll_main_dev12_inR42 = {main_dev1_in[99:0], 7'h2a};
  ZLL_Main_dev12  instR142 (zll_main_dev12_inR42[106:7], zll_main_dev12_inR42[6:0], zll_main_dev12_outR42);
  assign zll_main_dev12_inR43 = {main_dev1_in[99:0], 7'h2b};
  ZLL_Main_dev12  instR143 (zll_main_dev12_inR43[106:7], zll_main_dev12_inR43[6:0], zll_main_dev12_outR43);
  assign zll_main_dev12_inR44 = {main_dev1_in[99:0], 7'h2c};
  ZLL_Main_dev12  instR144 (zll_main_dev12_inR44[106:7], zll_main_dev12_inR44[6:0], zll_main_dev12_outR44);
  assign zll_main_dev12_inR45 = {main_dev1_in[99:0], 7'h2d};
  ZLL_Main_dev12  instR145 (zll_main_dev12_inR45[106:7], zll_main_dev12_inR45[6:0], zll_main_dev12_outR45);
  assign zll_main_dev12_inR46 = {main_dev1_in[99:0], 7'h2e};
  ZLL_Main_dev12  instR146 (zll_main_dev12_inR46[106:7], zll_main_dev12_inR46[6:0], zll_main_dev12_outR46);
  assign zll_main_dev12_inR47 = {main_dev1_in[99:0], 7'h2f};
  ZLL_Main_dev12  instR147 (zll_main_dev12_inR47[106:7], zll_main_dev12_inR47[6:0], zll_main_dev12_outR47);
  assign zll_main_dev12_inR48 = {main_dev1_in[99:0], 7'h30};
  ZLL_Main_dev12  instR148 (zll_main_dev12_inR48[106:7], zll_main_dev12_inR48[6:0], zll_main_dev12_outR48);
  assign zll_main_dev12_inR49 = {main_dev1_in[99:0], 7'h31};
  ZLL_Main_dev12  instR149 (zll_main_dev12_inR49[106:7], zll_main_dev12_inR49[6:0], zll_main_dev12_outR49);
  assign zll_main_dev12_inR50 = {main_dev1_in[99:0], 7'h32};
  ZLL_Main_dev12  instR150 (zll_main_dev12_inR50[106:7], zll_main_dev12_inR50[6:0], zll_main_dev12_outR50);
  assign zll_main_dev12_inR51 = {main_dev1_in[99:0], 7'h33};
  ZLL_Main_dev12  instR151 (zll_main_dev12_inR51[106:7], zll_main_dev12_inR51[6:0], zll_main_dev12_outR51);
  assign zll_main_dev12_inR52 = {main_dev1_in[99:0], 7'h34};
  ZLL_Main_dev12  instR152 (zll_main_dev12_inR52[106:7], zll_main_dev12_inR52[6:0], zll_main_dev12_outR52);
  assign zll_main_dev12_inR53 = {main_dev1_in[99:0], 7'h35};
  ZLL_Main_dev12  instR153 (zll_main_dev12_inR53[106:7], zll_main_dev12_inR53[6:0], zll_main_dev12_outR53);
  assign zll_main_dev12_inR54 = {main_dev1_in[99:0], 7'h36};
  ZLL_Main_dev12  instR154 (zll_main_dev12_inR54[106:7], zll_main_dev12_inR54[6:0], zll_main_dev12_outR54);
  assign zll_main_dev12_inR55 = {main_dev1_in[99:0], 7'h37};
  ZLL_Main_dev12  instR155 (zll_main_dev12_inR55[106:7], zll_main_dev12_inR55[6:0], zll_main_dev12_outR55);
  assign zll_main_dev12_inR56 = {main_dev1_in[99:0], 7'h38};
  ZLL_Main_dev12  instR156 (zll_main_dev12_inR56[106:7], zll_main_dev12_inR56[6:0], zll_main_dev12_outR56);
  assign zll_main_dev12_inR57 = {main_dev1_in[99:0], 7'h39};
  ZLL_Main_dev12  instR157 (zll_main_dev12_inR57[106:7], zll_main_dev12_inR57[6:0], zll_main_dev12_outR57);
  assign zll_main_dev12_inR58 = {main_dev1_in[99:0], 7'h3a};
  ZLL_Main_dev12  instR158 (zll_main_dev12_inR58[106:7], zll_main_dev12_inR58[6:0], zll_main_dev12_outR58);
  assign zll_main_dev12_inR59 = {main_dev1_in[99:0], 7'h3b};
  ZLL_Main_dev12  instR159 (zll_main_dev12_inR59[106:7], zll_main_dev12_inR59[6:0], zll_main_dev12_outR59);
  assign zll_main_dev12_inR60 = {main_dev1_in[99:0], 7'h3c};
  ZLL_Main_dev12  instR160 (zll_main_dev12_inR60[106:7], zll_main_dev12_inR60[6:0], zll_main_dev12_outR60);
  assign zll_main_dev12_inR61 = {main_dev1_in[99:0], 7'h3d};
  ZLL_Main_dev12  instR161 (zll_main_dev12_inR61[106:7], zll_main_dev12_inR61[6:0], zll_main_dev12_outR61);
  assign zll_main_dev12_inR62 = {main_dev1_in[99:0], 7'h3e};
  ZLL_Main_dev12  instR162 (zll_main_dev12_inR62[106:7], zll_main_dev12_inR62[6:0], zll_main_dev12_outR62);
  assign zll_main_dev12_inR63 = {main_dev1_in[99:0], 7'h3f};
  ZLL_Main_dev12  instR163 (zll_main_dev12_inR63[106:7], zll_main_dev12_inR63[6:0], zll_main_dev12_outR63);
  assign zll_main_dev12_inR64 = {main_dev1_in[99:0], 7'h40};
  ZLL_Main_dev12  instR164 (zll_main_dev12_inR64[106:7], zll_main_dev12_inR64[6:0], zll_main_dev12_outR64);
  assign zll_main_dev12_inR65 = {main_dev1_in[99:0], 7'h41};
  ZLL_Main_dev12  instR165 (zll_main_dev12_inR65[106:7], zll_main_dev12_inR65[6:0], zll_main_dev12_outR65);
  assign zll_main_dev12_inR66 = {main_dev1_in[99:0], 7'h42};
  ZLL_Main_dev12  instR166 (zll_main_dev12_inR66[106:7], zll_main_dev12_inR66[6:0], zll_main_dev12_outR66);
  assign zll_main_dev12_inR67 = {main_dev1_in[99:0], 7'h43};
  ZLL_Main_dev12  instR167 (zll_main_dev12_inR67[106:7], zll_main_dev12_inR67[6:0], zll_main_dev12_outR67);
  assign zll_main_dev12_inR68 = {main_dev1_in[99:0], 7'h44};
  ZLL_Main_dev12  instR168 (zll_main_dev12_inR68[106:7], zll_main_dev12_inR68[6:0], zll_main_dev12_outR68);
  assign zll_main_dev12_inR69 = {main_dev1_in[99:0], 7'h45};
  ZLL_Main_dev12  instR169 (zll_main_dev12_inR69[106:7], zll_main_dev12_inR69[6:0], zll_main_dev12_outR69);
  assign zll_main_dev12_inR70 = {main_dev1_in[99:0], 7'h46};
  ZLL_Main_dev12  instR170 (zll_main_dev12_inR70[106:7], zll_main_dev12_inR70[6:0], zll_main_dev12_outR70);
  assign zll_main_dev12_inR71 = {main_dev1_in[99:0], 7'h47};
  ZLL_Main_dev12  instR171 (zll_main_dev12_inR71[106:7], zll_main_dev12_inR71[6:0], zll_main_dev12_outR71);
  assign zll_main_dev12_inR72 = {main_dev1_in[99:0], 7'h48};
  ZLL_Main_dev12  instR172 (zll_main_dev12_inR72[106:7], zll_main_dev12_inR72[6:0], zll_main_dev12_outR72);
  assign zll_main_dev12_inR73 = {main_dev1_in[99:0], 7'h49};
  ZLL_Main_dev12  instR173 (zll_main_dev12_inR73[106:7], zll_main_dev12_inR73[6:0], zll_main_dev12_outR73);
  assign zll_main_dev12_inR74 = {main_dev1_in[99:0], 7'h4a};
  ZLL_Main_dev12  instR174 (zll_main_dev12_inR74[106:7], zll_main_dev12_inR74[6:0], zll_main_dev12_outR74);
  assign zll_main_dev12_inR75 = {main_dev1_in[99:0], 7'h4b};
  ZLL_Main_dev12  instR175 (zll_main_dev12_inR75[106:7], zll_main_dev12_inR75[6:0], zll_main_dev12_outR75);
  assign zll_main_dev12_inR76 = {main_dev1_in[99:0], 7'h4c};
  ZLL_Main_dev12  instR176 (zll_main_dev12_inR76[106:7], zll_main_dev12_inR76[6:0], zll_main_dev12_outR76);
  assign zll_main_dev12_inR77 = {main_dev1_in[99:0], 7'h4d};
  ZLL_Main_dev12  instR177 (zll_main_dev12_inR77[106:7], zll_main_dev12_inR77[6:0], zll_main_dev12_outR77);
  assign zll_main_dev12_inR78 = {main_dev1_in[99:0], 7'h4e};
  ZLL_Main_dev12  instR178 (zll_main_dev12_inR78[106:7], zll_main_dev12_inR78[6:0], zll_main_dev12_outR78);
  assign zll_main_dev12_inR79 = {main_dev1_in[99:0], 7'h4f};
  ZLL_Main_dev12  instR179 (zll_main_dev12_inR79[106:7], zll_main_dev12_inR79[6:0], zll_main_dev12_outR79);
  assign zll_main_dev12_inR80 = {main_dev1_in[99:0], 7'h50};
  ZLL_Main_dev12  instR180 (zll_main_dev12_inR80[106:7], zll_main_dev12_inR80[6:0], zll_main_dev12_outR80);
  assign zll_main_dev12_inR81 = {main_dev1_in[99:0], 7'h51};
  ZLL_Main_dev12  instR181 (zll_main_dev12_inR81[106:7], zll_main_dev12_inR81[6:0], zll_main_dev12_outR81);
  assign zll_main_dev12_inR82 = {main_dev1_in[99:0], 7'h52};
  ZLL_Main_dev12  instR182 (zll_main_dev12_inR82[106:7], zll_main_dev12_inR82[6:0], zll_main_dev12_outR82);
  assign zll_main_dev12_inR83 = {main_dev1_in[99:0], 7'h53};
  ZLL_Main_dev12  instR183 (zll_main_dev12_inR83[106:7], zll_main_dev12_inR83[6:0], zll_main_dev12_outR83);
  assign zll_main_dev12_inR84 = {main_dev1_in[99:0], 7'h54};
  ZLL_Main_dev12  instR184 (zll_main_dev12_inR84[106:7], zll_main_dev12_inR84[6:0], zll_main_dev12_outR84);
  assign zll_main_dev12_inR85 = {main_dev1_in[99:0], 7'h55};
  ZLL_Main_dev12  instR185 (zll_main_dev12_inR85[106:7], zll_main_dev12_inR85[6:0], zll_main_dev12_outR85);
  assign zll_main_dev12_inR86 = {main_dev1_in[99:0], 7'h56};
  ZLL_Main_dev12  instR186 (zll_main_dev12_inR86[106:7], zll_main_dev12_inR86[6:0], zll_main_dev12_outR86);
  assign zll_main_dev12_inR87 = {main_dev1_in[99:0], 7'h57};
  ZLL_Main_dev12  instR187 (zll_main_dev12_inR87[106:7], zll_main_dev12_inR87[6:0], zll_main_dev12_outR87);
  assign zll_main_dev12_inR88 = {main_dev1_in[99:0], 7'h58};
  ZLL_Main_dev12  instR188 (zll_main_dev12_inR88[106:7], zll_main_dev12_inR88[6:0], zll_main_dev12_outR88);
  assign zll_main_dev12_inR89 = {main_dev1_in[99:0], 7'h59};
  ZLL_Main_dev12  instR189 (zll_main_dev12_inR89[106:7], zll_main_dev12_inR89[6:0], zll_main_dev12_outR89);
  assign zll_main_dev12_inR90 = {main_dev1_in[99:0], 7'h5a};
  ZLL_Main_dev12  instR190 (zll_main_dev12_inR90[106:7], zll_main_dev12_inR90[6:0], zll_main_dev12_outR90);
  assign zll_main_dev12_inR91 = {main_dev1_in[99:0], 7'h5b};
  ZLL_Main_dev12  instR191 (zll_main_dev12_inR91[106:7], zll_main_dev12_inR91[6:0], zll_main_dev12_outR91);
  assign zll_main_dev12_inR92 = {main_dev1_in[99:0], 7'h5c};
  ZLL_Main_dev12  instR192 (zll_main_dev12_inR92[106:7], zll_main_dev12_inR92[6:0], zll_main_dev12_outR92);
  assign zll_main_dev12_inR93 = {main_dev1_in[99:0], 7'h5d};
  ZLL_Main_dev12  instR193 (zll_main_dev12_inR93[106:7], zll_main_dev12_inR93[6:0], zll_main_dev12_outR93);
  assign zll_main_dev12_inR94 = {main_dev1_in[99:0], 7'h5e};
  ZLL_Main_dev12  instR194 (zll_main_dev12_inR94[106:7], zll_main_dev12_inR94[6:0], zll_main_dev12_outR94);
  assign zll_main_dev12_inR95 = {main_dev1_in[99:0], 7'h5f};
  ZLL_Main_dev12  instR195 (zll_main_dev12_inR95[106:7], zll_main_dev12_inR95[6:0], zll_main_dev12_outR95);
  assign zll_main_dev12_inR96 = {main_dev1_in[99:0], 7'h60};
  ZLL_Main_dev12  instR196 (zll_main_dev12_inR96[106:7], zll_main_dev12_inR96[6:0], zll_main_dev12_outR96);
  assign zll_main_dev12_inR97 = {main_dev1_in[99:0], 7'h61};
  ZLL_Main_dev12  instR197 (zll_main_dev12_inR97[106:7], zll_main_dev12_inR97[6:0], zll_main_dev12_outR97);
  assign zll_main_dev12_inR98 = {main_dev1_in[99:0], 7'h62};
  ZLL_Main_dev12  instR198 (zll_main_dev12_inR98[106:7], zll_main_dev12_inR98[6:0], zll_main_dev12_outR98);
  assign zll_main_dev12_inR99 = {main_dev1_in[99:0], 7'h63};
  ZLL_Main_dev12  instR199 (zll_main_dev12_inR99[106:7], zll_main_dev12_inR99[6:0], zll_main_dev12_outR99);
  assign zll_main_dev15_in = {main_dev1_in[99:0], 7'h0};
  ZLL_Main_dev15  instR200 (zll_main_dev15_in[106:7], zll_main_dev15_in[6:0], zll_main_dev15_out);
  assign zll_main_dev15_inR1 = {main_dev1_in[99:0], 7'h1};
  ZLL_Main_dev15  instR201 (zll_main_dev15_inR1[106:7], zll_main_dev15_inR1[6:0], zll_main_dev15_outR1);
  assign zll_main_dev15_inR2 = {main_dev1_in[99:0], 7'h2};
  ZLL_Main_dev15  instR202 (zll_main_dev15_inR2[106:7], zll_main_dev15_inR2[6:0], zll_main_dev15_outR2);
  assign zll_main_dev15_inR3 = {main_dev1_in[99:0], 7'h3};
  ZLL_Main_dev15  instR203 (zll_main_dev15_inR3[106:7], zll_main_dev15_inR3[6:0], zll_main_dev15_outR3);
  assign zll_main_dev15_inR4 = {main_dev1_in[99:0], 7'h4};
  ZLL_Main_dev15  instR204 (zll_main_dev15_inR4[106:7], zll_main_dev15_inR4[6:0], zll_main_dev15_outR4);
  assign zll_main_dev15_inR5 = {main_dev1_in[99:0], 7'h5};
  ZLL_Main_dev15  instR205 (zll_main_dev15_inR5[106:7], zll_main_dev15_inR5[6:0], zll_main_dev15_outR5);
  assign zll_main_dev15_inR6 = {main_dev1_in[99:0], 7'h6};
  ZLL_Main_dev15  instR206 (zll_main_dev15_inR6[106:7], zll_main_dev15_inR6[6:0], zll_main_dev15_outR6);
  assign zll_main_dev15_inR7 = {main_dev1_in[99:0], 7'h7};
  ZLL_Main_dev15  instR207 (zll_main_dev15_inR7[106:7], zll_main_dev15_inR7[6:0], zll_main_dev15_outR7);
  assign zll_main_dev15_inR8 = {main_dev1_in[99:0], 7'h8};
  ZLL_Main_dev15  instR208 (zll_main_dev15_inR8[106:7], zll_main_dev15_inR8[6:0], zll_main_dev15_outR8);
  assign zll_main_dev15_inR9 = {main_dev1_in[99:0], 7'h9};
  ZLL_Main_dev15  instR209 (zll_main_dev15_inR9[106:7], zll_main_dev15_inR9[6:0], zll_main_dev15_outR9);
  assign zll_main_dev15_inR10 = {main_dev1_in[99:0], 7'ha};
  ZLL_Main_dev15  instR210 (zll_main_dev15_inR10[106:7], zll_main_dev15_inR10[6:0], zll_main_dev15_outR10);
  assign zll_main_dev15_inR11 = {main_dev1_in[99:0], 7'hb};
  ZLL_Main_dev15  instR211 (zll_main_dev15_inR11[106:7], zll_main_dev15_inR11[6:0], zll_main_dev15_outR11);
  assign zll_main_dev15_inR12 = {main_dev1_in[99:0], 7'hc};
  ZLL_Main_dev15  instR212 (zll_main_dev15_inR12[106:7], zll_main_dev15_inR12[6:0], zll_main_dev15_outR12);
  assign zll_main_dev15_inR13 = {main_dev1_in[99:0], 7'hd};
  ZLL_Main_dev15  instR213 (zll_main_dev15_inR13[106:7], zll_main_dev15_inR13[6:0], zll_main_dev15_outR13);
  assign zll_main_dev15_inR14 = {main_dev1_in[99:0], 7'he};
  ZLL_Main_dev15  instR214 (zll_main_dev15_inR14[106:7], zll_main_dev15_inR14[6:0], zll_main_dev15_outR14);
  assign zll_main_dev15_inR15 = {main_dev1_in[99:0], 7'hf};
  ZLL_Main_dev15  instR215 (zll_main_dev15_inR15[106:7], zll_main_dev15_inR15[6:0], zll_main_dev15_outR15);
  assign zll_main_dev15_inR16 = {main_dev1_in[99:0], 7'h10};
  ZLL_Main_dev15  instR216 (zll_main_dev15_inR16[106:7], zll_main_dev15_inR16[6:0], zll_main_dev15_outR16);
  assign zll_main_dev15_inR17 = {main_dev1_in[99:0], 7'h11};
  ZLL_Main_dev15  instR217 (zll_main_dev15_inR17[106:7], zll_main_dev15_inR17[6:0], zll_main_dev15_outR17);
  assign zll_main_dev15_inR18 = {main_dev1_in[99:0], 7'h12};
  ZLL_Main_dev15  instR218 (zll_main_dev15_inR18[106:7], zll_main_dev15_inR18[6:0], zll_main_dev15_outR18);
  assign zll_main_dev15_inR19 = {main_dev1_in[99:0], 7'h13};
  ZLL_Main_dev15  instR219 (zll_main_dev15_inR19[106:7], zll_main_dev15_inR19[6:0], zll_main_dev15_outR19);
  assign zll_main_dev15_inR20 = {main_dev1_in[99:0], 7'h14};
  ZLL_Main_dev15  instR220 (zll_main_dev15_inR20[106:7], zll_main_dev15_inR20[6:0], zll_main_dev15_outR20);
  assign zll_main_dev15_inR21 = {main_dev1_in[99:0], 7'h15};
  ZLL_Main_dev15  instR221 (zll_main_dev15_inR21[106:7], zll_main_dev15_inR21[6:0], zll_main_dev15_outR21);
  assign zll_main_dev15_inR22 = {main_dev1_in[99:0], 7'h16};
  ZLL_Main_dev15  instR222 (zll_main_dev15_inR22[106:7], zll_main_dev15_inR22[6:0], zll_main_dev15_outR22);
  assign zll_main_dev15_inR23 = {main_dev1_in[99:0], 7'h17};
  ZLL_Main_dev15  instR223 (zll_main_dev15_inR23[106:7], zll_main_dev15_inR23[6:0], zll_main_dev15_outR23);
  assign zll_main_dev15_inR24 = {main_dev1_in[99:0], 7'h18};
  ZLL_Main_dev15  instR224 (zll_main_dev15_inR24[106:7], zll_main_dev15_inR24[6:0], zll_main_dev15_outR24);
  assign zll_main_dev15_inR25 = {main_dev1_in[99:0], 7'h19};
  ZLL_Main_dev15  instR225 (zll_main_dev15_inR25[106:7], zll_main_dev15_inR25[6:0], zll_main_dev15_outR25);
  assign zll_main_dev15_inR26 = {main_dev1_in[99:0], 7'h1a};
  ZLL_Main_dev15  instR226 (zll_main_dev15_inR26[106:7], zll_main_dev15_inR26[6:0], zll_main_dev15_outR26);
  assign zll_main_dev15_inR27 = {main_dev1_in[99:0], 7'h1b};
  ZLL_Main_dev15  instR227 (zll_main_dev15_inR27[106:7], zll_main_dev15_inR27[6:0], zll_main_dev15_outR27);
  assign zll_main_dev15_inR28 = {main_dev1_in[99:0], 7'h1c};
  ZLL_Main_dev15  instR228 (zll_main_dev15_inR28[106:7], zll_main_dev15_inR28[6:0], zll_main_dev15_outR28);
  assign zll_main_dev15_inR29 = {main_dev1_in[99:0], 7'h1d};
  ZLL_Main_dev15  instR229 (zll_main_dev15_inR29[106:7], zll_main_dev15_inR29[6:0], zll_main_dev15_outR29);
  assign zll_main_dev15_inR30 = {main_dev1_in[99:0], 7'h1e};
  ZLL_Main_dev15  instR230 (zll_main_dev15_inR30[106:7], zll_main_dev15_inR30[6:0], zll_main_dev15_outR30);
  assign zll_main_dev15_inR31 = {main_dev1_in[99:0], 7'h1f};
  ZLL_Main_dev15  instR231 (zll_main_dev15_inR31[106:7], zll_main_dev15_inR31[6:0], zll_main_dev15_outR31);
  assign zll_main_dev15_inR32 = {main_dev1_in[99:0], 7'h20};
  ZLL_Main_dev15  instR232 (zll_main_dev15_inR32[106:7], zll_main_dev15_inR32[6:0], zll_main_dev15_outR32);
  assign zll_main_dev15_inR33 = {main_dev1_in[99:0], 7'h21};
  ZLL_Main_dev15  instR233 (zll_main_dev15_inR33[106:7], zll_main_dev15_inR33[6:0], zll_main_dev15_outR33);
  assign zll_main_dev15_inR34 = {main_dev1_in[99:0], 7'h22};
  ZLL_Main_dev15  instR234 (zll_main_dev15_inR34[106:7], zll_main_dev15_inR34[6:0], zll_main_dev15_outR34);
  assign zll_main_dev15_inR35 = {main_dev1_in[99:0], 7'h23};
  ZLL_Main_dev15  instR235 (zll_main_dev15_inR35[106:7], zll_main_dev15_inR35[6:0], zll_main_dev15_outR35);
  assign zll_main_dev15_inR36 = {main_dev1_in[99:0], 7'h24};
  ZLL_Main_dev15  instR236 (zll_main_dev15_inR36[106:7], zll_main_dev15_inR36[6:0], zll_main_dev15_outR36);
  assign zll_main_dev15_inR37 = {main_dev1_in[99:0], 7'h25};
  ZLL_Main_dev15  instR237 (zll_main_dev15_inR37[106:7], zll_main_dev15_inR37[6:0], zll_main_dev15_outR37);
  assign zll_main_dev15_inR38 = {main_dev1_in[99:0], 7'h26};
  ZLL_Main_dev15  instR238 (zll_main_dev15_inR38[106:7], zll_main_dev15_inR38[6:0], zll_main_dev15_outR38);
  assign zll_main_dev15_inR39 = {main_dev1_in[99:0], 7'h27};
  ZLL_Main_dev15  instR239 (zll_main_dev15_inR39[106:7], zll_main_dev15_inR39[6:0], zll_main_dev15_outR39);
  assign zll_main_dev15_inR40 = {main_dev1_in[99:0], 7'h28};
  ZLL_Main_dev15  instR240 (zll_main_dev15_inR40[106:7], zll_main_dev15_inR40[6:0], zll_main_dev15_outR40);
  assign zll_main_dev15_inR41 = {main_dev1_in[99:0], 7'h29};
  ZLL_Main_dev15  instR241 (zll_main_dev15_inR41[106:7], zll_main_dev15_inR41[6:0], zll_main_dev15_outR41);
  assign zll_main_dev15_inR42 = {main_dev1_in[99:0], 7'h2a};
  ZLL_Main_dev15  instR242 (zll_main_dev15_inR42[106:7], zll_main_dev15_inR42[6:0], zll_main_dev15_outR42);
  assign zll_main_dev15_inR43 = {main_dev1_in[99:0], 7'h2b};
  ZLL_Main_dev15  instR243 (zll_main_dev15_inR43[106:7], zll_main_dev15_inR43[6:0], zll_main_dev15_outR43);
  assign zll_main_dev15_inR44 = {main_dev1_in[99:0], 7'h2c};
  ZLL_Main_dev15  instR244 (zll_main_dev15_inR44[106:7], zll_main_dev15_inR44[6:0], zll_main_dev15_outR44);
  assign zll_main_dev15_inR45 = {main_dev1_in[99:0], 7'h2d};
  ZLL_Main_dev15  instR245 (zll_main_dev15_inR45[106:7], zll_main_dev15_inR45[6:0], zll_main_dev15_outR45);
  assign zll_main_dev15_inR46 = {main_dev1_in[99:0], 7'h2e};
  ZLL_Main_dev15  instR246 (zll_main_dev15_inR46[106:7], zll_main_dev15_inR46[6:0], zll_main_dev15_outR46);
  assign zll_main_dev15_inR47 = {main_dev1_in[99:0], 7'h2f};
  ZLL_Main_dev15  instR247 (zll_main_dev15_inR47[106:7], zll_main_dev15_inR47[6:0], zll_main_dev15_outR47);
  assign zll_main_dev15_inR48 = {main_dev1_in[99:0], 7'h30};
  ZLL_Main_dev15  instR248 (zll_main_dev15_inR48[106:7], zll_main_dev15_inR48[6:0], zll_main_dev15_outR48);
  assign zll_main_dev15_inR49 = {main_dev1_in[99:0], 7'h31};
  ZLL_Main_dev15  instR249 (zll_main_dev15_inR49[106:7], zll_main_dev15_inR49[6:0], zll_main_dev15_outR49);
  assign zll_main_dev15_inR50 = {main_dev1_in[99:0], 7'h32};
  ZLL_Main_dev15  instR250 (zll_main_dev15_inR50[106:7], zll_main_dev15_inR50[6:0], zll_main_dev15_outR50);
  assign zll_main_dev15_inR51 = {main_dev1_in[99:0], 7'h33};
  ZLL_Main_dev15  instR251 (zll_main_dev15_inR51[106:7], zll_main_dev15_inR51[6:0], zll_main_dev15_outR51);
  assign zll_main_dev15_inR52 = {main_dev1_in[99:0], 7'h34};
  ZLL_Main_dev15  instR252 (zll_main_dev15_inR52[106:7], zll_main_dev15_inR52[6:0], zll_main_dev15_outR52);
  assign zll_main_dev15_inR53 = {main_dev1_in[99:0], 7'h35};
  ZLL_Main_dev15  instR253 (zll_main_dev15_inR53[106:7], zll_main_dev15_inR53[6:0], zll_main_dev15_outR53);
  assign zll_main_dev15_inR54 = {main_dev1_in[99:0], 7'h36};
  ZLL_Main_dev15  instR254 (zll_main_dev15_inR54[106:7], zll_main_dev15_inR54[6:0], zll_main_dev15_outR54);
  assign zll_main_dev15_inR55 = {main_dev1_in[99:0], 7'h37};
  ZLL_Main_dev15  instR255 (zll_main_dev15_inR55[106:7], zll_main_dev15_inR55[6:0], zll_main_dev15_outR55);
  assign zll_main_dev15_inR56 = {main_dev1_in[99:0], 7'h38};
  ZLL_Main_dev15  instR256 (zll_main_dev15_inR56[106:7], zll_main_dev15_inR56[6:0], zll_main_dev15_outR56);
  assign zll_main_dev15_inR57 = {main_dev1_in[99:0], 7'h39};
  ZLL_Main_dev15  instR257 (zll_main_dev15_inR57[106:7], zll_main_dev15_inR57[6:0], zll_main_dev15_outR57);
  assign zll_main_dev15_inR58 = {main_dev1_in[99:0], 7'h3a};
  ZLL_Main_dev15  instR258 (zll_main_dev15_inR58[106:7], zll_main_dev15_inR58[6:0], zll_main_dev15_outR58);
  assign zll_main_dev15_inR59 = {main_dev1_in[99:0], 7'h3b};
  ZLL_Main_dev15  instR259 (zll_main_dev15_inR59[106:7], zll_main_dev15_inR59[6:0], zll_main_dev15_outR59);
  assign zll_main_dev15_inR60 = {main_dev1_in[99:0], 7'h3c};
  ZLL_Main_dev15  instR260 (zll_main_dev15_inR60[106:7], zll_main_dev15_inR60[6:0], zll_main_dev15_outR60);
  assign zll_main_dev15_inR61 = {main_dev1_in[99:0], 7'h3d};
  ZLL_Main_dev15  instR261 (zll_main_dev15_inR61[106:7], zll_main_dev15_inR61[6:0], zll_main_dev15_outR61);
  assign zll_main_dev15_inR62 = {main_dev1_in[99:0], 7'h3e};
  ZLL_Main_dev15  instR262 (zll_main_dev15_inR62[106:7], zll_main_dev15_inR62[6:0], zll_main_dev15_outR62);
  assign zll_main_dev15_inR63 = {main_dev1_in[99:0], 7'h3f};
  ZLL_Main_dev15  instR263 (zll_main_dev15_inR63[106:7], zll_main_dev15_inR63[6:0], zll_main_dev15_outR63);
  assign zll_main_dev15_inR64 = {main_dev1_in[99:0], 7'h40};
  ZLL_Main_dev15  instR264 (zll_main_dev15_inR64[106:7], zll_main_dev15_inR64[6:0], zll_main_dev15_outR64);
  assign zll_main_dev15_inR65 = {main_dev1_in[99:0], 7'h41};
  ZLL_Main_dev15  instR265 (zll_main_dev15_inR65[106:7], zll_main_dev15_inR65[6:0], zll_main_dev15_outR65);
  assign zll_main_dev15_inR66 = {main_dev1_in[99:0], 7'h42};
  ZLL_Main_dev15  instR266 (zll_main_dev15_inR66[106:7], zll_main_dev15_inR66[6:0], zll_main_dev15_outR66);
  assign zll_main_dev15_inR67 = {main_dev1_in[99:0], 7'h43};
  ZLL_Main_dev15  instR267 (zll_main_dev15_inR67[106:7], zll_main_dev15_inR67[6:0], zll_main_dev15_outR67);
  assign zll_main_dev15_inR68 = {main_dev1_in[99:0], 7'h44};
  ZLL_Main_dev15  instR268 (zll_main_dev15_inR68[106:7], zll_main_dev15_inR68[6:0], zll_main_dev15_outR68);
  assign zll_main_dev15_inR69 = {main_dev1_in[99:0], 7'h45};
  ZLL_Main_dev15  instR269 (zll_main_dev15_inR69[106:7], zll_main_dev15_inR69[6:0], zll_main_dev15_outR69);
  assign zll_main_dev15_inR70 = {main_dev1_in[99:0], 7'h46};
  ZLL_Main_dev15  instR270 (zll_main_dev15_inR70[106:7], zll_main_dev15_inR70[6:0], zll_main_dev15_outR70);
  assign zll_main_dev15_inR71 = {main_dev1_in[99:0], 7'h47};
  ZLL_Main_dev15  instR271 (zll_main_dev15_inR71[106:7], zll_main_dev15_inR71[6:0], zll_main_dev15_outR71);
  assign zll_main_dev15_inR72 = {main_dev1_in[99:0], 7'h48};
  ZLL_Main_dev15  instR272 (zll_main_dev15_inR72[106:7], zll_main_dev15_inR72[6:0], zll_main_dev15_outR72);
  assign zll_main_dev15_inR73 = {main_dev1_in[99:0], 7'h49};
  ZLL_Main_dev15  instR273 (zll_main_dev15_inR73[106:7], zll_main_dev15_inR73[6:0], zll_main_dev15_outR73);
  assign zll_main_dev15_inR74 = {main_dev1_in[99:0], 7'h4a};
  ZLL_Main_dev15  instR274 (zll_main_dev15_inR74[106:7], zll_main_dev15_inR74[6:0], zll_main_dev15_outR74);
  assign zll_main_dev15_inR75 = {main_dev1_in[99:0], 7'h4b};
  ZLL_Main_dev15  instR275 (zll_main_dev15_inR75[106:7], zll_main_dev15_inR75[6:0], zll_main_dev15_outR75);
  assign zll_main_dev15_inR76 = {main_dev1_in[99:0], 7'h4c};
  ZLL_Main_dev15  instR276 (zll_main_dev15_inR76[106:7], zll_main_dev15_inR76[6:0], zll_main_dev15_outR76);
  assign zll_main_dev15_inR77 = {main_dev1_in[99:0], 7'h4d};
  ZLL_Main_dev15  instR277 (zll_main_dev15_inR77[106:7], zll_main_dev15_inR77[6:0], zll_main_dev15_outR77);
  assign zll_main_dev15_inR78 = {main_dev1_in[99:0], 7'h4e};
  ZLL_Main_dev15  instR278 (zll_main_dev15_inR78[106:7], zll_main_dev15_inR78[6:0], zll_main_dev15_outR78);
  assign zll_main_dev15_inR79 = {main_dev1_in[99:0], 7'h4f};
  ZLL_Main_dev15  instR279 (zll_main_dev15_inR79[106:7], zll_main_dev15_inR79[6:0], zll_main_dev15_outR79);
  assign zll_main_dev15_inR80 = {main_dev1_in[99:0], 7'h50};
  ZLL_Main_dev15  instR280 (zll_main_dev15_inR80[106:7], zll_main_dev15_inR80[6:0], zll_main_dev15_outR80);
  assign zll_main_dev15_inR81 = {main_dev1_in[99:0], 7'h51};
  ZLL_Main_dev15  instR281 (zll_main_dev15_inR81[106:7], zll_main_dev15_inR81[6:0], zll_main_dev15_outR81);
  assign zll_main_dev15_inR82 = {main_dev1_in[99:0], 7'h52};
  ZLL_Main_dev15  instR282 (zll_main_dev15_inR82[106:7], zll_main_dev15_inR82[6:0], zll_main_dev15_outR82);
  assign zll_main_dev15_inR83 = {main_dev1_in[99:0], 7'h53};
  ZLL_Main_dev15  instR283 (zll_main_dev15_inR83[106:7], zll_main_dev15_inR83[6:0], zll_main_dev15_outR83);
  assign zll_main_dev15_inR84 = {main_dev1_in[99:0], 7'h54};
  ZLL_Main_dev15  instR284 (zll_main_dev15_inR84[106:7], zll_main_dev15_inR84[6:0], zll_main_dev15_outR84);
  assign zll_main_dev15_inR85 = {main_dev1_in[99:0], 7'h55};
  ZLL_Main_dev15  instR285 (zll_main_dev15_inR85[106:7], zll_main_dev15_inR85[6:0], zll_main_dev15_outR85);
  assign zll_main_dev15_inR86 = {main_dev1_in[99:0], 7'h56};
  ZLL_Main_dev15  instR286 (zll_main_dev15_inR86[106:7], zll_main_dev15_inR86[6:0], zll_main_dev15_outR86);
  assign zll_main_dev15_inR87 = {main_dev1_in[99:0], 7'h57};
  ZLL_Main_dev15  instR287 (zll_main_dev15_inR87[106:7], zll_main_dev15_inR87[6:0], zll_main_dev15_outR87);
  assign zll_main_dev15_inR88 = {main_dev1_in[99:0], 7'h58};
  ZLL_Main_dev15  instR288 (zll_main_dev15_inR88[106:7], zll_main_dev15_inR88[6:0], zll_main_dev15_outR88);
  assign zll_main_dev15_inR89 = {main_dev1_in[99:0], 7'h59};
  ZLL_Main_dev15  instR289 (zll_main_dev15_inR89[106:7], zll_main_dev15_inR89[6:0], zll_main_dev15_outR89);
  assign zll_main_dev15_inR90 = {main_dev1_in[99:0], 7'h5a};
  ZLL_Main_dev15  instR290 (zll_main_dev15_inR90[106:7], zll_main_dev15_inR90[6:0], zll_main_dev15_outR90);
  assign zll_main_dev15_inR91 = {main_dev1_in[99:0], 7'h5b};
  ZLL_Main_dev15  instR291 (zll_main_dev15_inR91[106:7], zll_main_dev15_inR91[6:0], zll_main_dev15_outR91);
  assign zll_main_dev15_inR92 = {main_dev1_in[99:0], 7'h5c};
  ZLL_Main_dev15  instR292 (zll_main_dev15_inR92[106:7], zll_main_dev15_inR92[6:0], zll_main_dev15_outR92);
  assign zll_main_dev15_inR93 = {main_dev1_in[99:0], 7'h5d};
  ZLL_Main_dev15  instR293 (zll_main_dev15_inR93[106:7], zll_main_dev15_inR93[6:0], zll_main_dev15_outR93);
  assign zll_main_dev15_inR94 = {main_dev1_in[99:0], 7'h5e};
  ZLL_Main_dev15  instR294 (zll_main_dev15_inR94[106:7], zll_main_dev15_inR94[6:0], zll_main_dev15_outR94);
  assign zll_main_dev15_inR95 = {main_dev1_in[99:0], 7'h5f};
  ZLL_Main_dev15  instR295 (zll_main_dev15_inR95[106:7], zll_main_dev15_inR95[6:0], zll_main_dev15_outR95);
  assign zll_main_dev15_inR96 = {main_dev1_in[99:0], 7'h60};
  ZLL_Main_dev15  instR296 (zll_main_dev15_inR96[106:7], zll_main_dev15_inR96[6:0], zll_main_dev15_outR96);
  assign zll_main_dev15_inR97 = {main_dev1_in[99:0], 7'h61};
  ZLL_Main_dev15  instR297 (zll_main_dev15_inR97[106:7], zll_main_dev15_inR97[6:0], zll_main_dev15_outR97);
  assign zll_main_dev15_inR98 = {main_dev1_in[99:0], 7'h62};
  ZLL_Main_dev15  instR298 (zll_main_dev15_inR98[106:7], zll_main_dev15_inR98[6:0], zll_main_dev15_outR98);
  assign zll_main_dev15_inR99 = {main_dev1_in[99:0], 7'h63};
  ZLL_Main_dev15  instR299 (zll_main_dev15_inR99[106:7], zll_main_dev15_inR99[6:0], zll_main_dev15_outR99);
  assign zll_main_dev8_in = {main_dev1_in[99:0], 7'h0};
  ZLL_Main_dev8  instR300 (zll_main_dev8_in[106:7], zll_main_dev8_in[6:0], zll_main_dev8_out);
  assign zll_main_dev8_inR1 = {main_dev1_in[99:0], 7'h1};
  ZLL_Main_dev8  instR301 (zll_main_dev8_inR1[106:7], zll_main_dev8_inR1[6:0], zll_main_dev8_outR1);
  assign zll_main_dev8_inR2 = {main_dev1_in[99:0], 7'h2};
  ZLL_Main_dev8  instR302 (zll_main_dev8_inR2[106:7], zll_main_dev8_inR2[6:0], zll_main_dev8_outR2);
  assign zll_main_dev8_inR3 = {main_dev1_in[99:0], 7'h3};
  ZLL_Main_dev8  instR303 (zll_main_dev8_inR3[106:7], zll_main_dev8_inR3[6:0], zll_main_dev8_outR3);
  assign zll_main_dev8_inR4 = {main_dev1_in[99:0], 7'h4};
  ZLL_Main_dev8  instR304 (zll_main_dev8_inR4[106:7], zll_main_dev8_inR4[6:0], zll_main_dev8_outR4);
  assign zll_main_dev8_inR5 = {main_dev1_in[99:0], 7'h5};
  ZLL_Main_dev8  instR305 (zll_main_dev8_inR5[106:7], zll_main_dev8_inR5[6:0], zll_main_dev8_outR5);
  assign zll_main_dev8_inR6 = {main_dev1_in[99:0], 7'h6};
  ZLL_Main_dev8  instR306 (zll_main_dev8_inR6[106:7], zll_main_dev8_inR6[6:0], zll_main_dev8_outR6);
  assign zll_main_dev8_inR7 = {main_dev1_in[99:0], 7'h7};
  ZLL_Main_dev8  instR307 (zll_main_dev8_inR7[106:7], zll_main_dev8_inR7[6:0], zll_main_dev8_outR7);
  assign zll_main_dev8_inR8 = {main_dev1_in[99:0], 7'h8};
  ZLL_Main_dev8  instR308 (zll_main_dev8_inR8[106:7], zll_main_dev8_inR8[6:0], zll_main_dev8_outR8);
  assign zll_main_dev8_inR9 = {main_dev1_in[99:0], 7'h9};
  ZLL_Main_dev8  instR309 (zll_main_dev8_inR9[106:7], zll_main_dev8_inR9[6:0], zll_main_dev8_outR9);
  assign zll_main_dev8_inR10 = {main_dev1_in[99:0], 7'ha};
  ZLL_Main_dev8  instR310 (zll_main_dev8_inR10[106:7], zll_main_dev8_inR10[6:0], zll_main_dev8_outR10);
  assign zll_main_dev8_inR11 = {main_dev1_in[99:0], 7'hb};
  ZLL_Main_dev8  instR311 (zll_main_dev8_inR11[106:7], zll_main_dev8_inR11[6:0], zll_main_dev8_outR11);
  assign zll_main_dev8_inR12 = {main_dev1_in[99:0], 7'hc};
  ZLL_Main_dev8  instR312 (zll_main_dev8_inR12[106:7], zll_main_dev8_inR12[6:0], zll_main_dev8_outR12);
  assign zll_main_dev8_inR13 = {main_dev1_in[99:0], 7'hd};
  ZLL_Main_dev8  instR313 (zll_main_dev8_inR13[106:7], zll_main_dev8_inR13[6:0], zll_main_dev8_outR13);
  assign zll_main_dev8_inR14 = {main_dev1_in[99:0], 7'he};
  ZLL_Main_dev8  instR314 (zll_main_dev8_inR14[106:7], zll_main_dev8_inR14[6:0], zll_main_dev8_outR14);
  assign zll_main_dev8_inR15 = {main_dev1_in[99:0], 7'hf};
  ZLL_Main_dev8  instR315 (zll_main_dev8_inR15[106:7], zll_main_dev8_inR15[6:0], zll_main_dev8_outR15);
  assign zll_main_dev8_inR16 = {main_dev1_in[99:0], 7'h10};
  ZLL_Main_dev8  instR316 (zll_main_dev8_inR16[106:7], zll_main_dev8_inR16[6:0], zll_main_dev8_outR16);
  assign zll_main_dev8_inR17 = {main_dev1_in[99:0], 7'h11};
  ZLL_Main_dev8  instR317 (zll_main_dev8_inR17[106:7], zll_main_dev8_inR17[6:0], zll_main_dev8_outR17);
  assign zll_main_dev8_inR18 = {main_dev1_in[99:0], 7'h12};
  ZLL_Main_dev8  instR318 (zll_main_dev8_inR18[106:7], zll_main_dev8_inR18[6:0], zll_main_dev8_outR18);
  assign zll_main_dev8_inR19 = {main_dev1_in[99:0], 7'h13};
  ZLL_Main_dev8  instR319 (zll_main_dev8_inR19[106:7], zll_main_dev8_inR19[6:0], zll_main_dev8_outR19);
  assign zll_main_dev8_inR20 = {main_dev1_in[99:0], 7'h14};
  ZLL_Main_dev8  instR320 (zll_main_dev8_inR20[106:7], zll_main_dev8_inR20[6:0], zll_main_dev8_outR20);
  assign zll_main_dev8_inR21 = {main_dev1_in[99:0], 7'h15};
  ZLL_Main_dev8  instR321 (zll_main_dev8_inR21[106:7], zll_main_dev8_inR21[6:0], zll_main_dev8_outR21);
  assign zll_main_dev8_inR22 = {main_dev1_in[99:0], 7'h16};
  ZLL_Main_dev8  instR322 (zll_main_dev8_inR22[106:7], zll_main_dev8_inR22[6:0], zll_main_dev8_outR22);
  assign zll_main_dev8_inR23 = {main_dev1_in[99:0], 7'h17};
  ZLL_Main_dev8  instR323 (zll_main_dev8_inR23[106:7], zll_main_dev8_inR23[6:0], zll_main_dev8_outR23);
  assign zll_main_dev8_inR24 = {main_dev1_in[99:0], 7'h18};
  ZLL_Main_dev8  instR324 (zll_main_dev8_inR24[106:7], zll_main_dev8_inR24[6:0], zll_main_dev8_outR24);
  assign zll_main_dev8_inR25 = {main_dev1_in[99:0], 7'h19};
  ZLL_Main_dev8  instR325 (zll_main_dev8_inR25[106:7], zll_main_dev8_inR25[6:0], zll_main_dev8_outR25);
  assign zll_main_dev8_inR26 = {main_dev1_in[99:0], 7'h1a};
  ZLL_Main_dev8  instR326 (zll_main_dev8_inR26[106:7], zll_main_dev8_inR26[6:0], zll_main_dev8_outR26);
  assign zll_main_dev8_inR27 = {main_dev1_in[99:0], 7'h1b};
  ZLL_Main_dev8  instR327 (zll_main_dev8_inR27[106:7], zll_main_dev8_inR27[6:0], zll_main_dev8_outR27);
  assign zll_main_dev8_inR28 = {main_dev1_in[99:0], 7'h1c};
  ZLL_Main_dev8  instR328 (zll_main_dev8_inR28[106:7], zll_main_dev8_inR28[6:0], zll_main_dev8_outR28);
  assign zll_main_dev8_inR29 = {main_dev1_in[99:0], 7'h1d};
  ZLL_Main_dev8  instR329 (zll_main_dev8_inR29[106:7], zll_main_dev8_inR29[6:0], zll_main_dev8_outR29);
  assign zll_main_dev8_inR30 = {main_dev1_in[99:0], 7'h1e};
  ZLL_Main_dev8  instR330 (zll_main_dev8_inR30[106:7], zll_main_dev8_inR30[6:0], zll_main_dev8_outR30);
  assign zll_main_dev8_inR31 = {main_dev1_in[99:0], 7'h1f};
  ZLL_Main_dev8  instR331 (zll_main_dev8_inR31[106:7], zll_main_dev8_inR31[6:0], zll_main_dev8_outR31);
  assign zll_main_dev8_inR32 = {main_dev1_in[99:0], 7'h20};
  ZLL_Main_dev8  instR332 (zll_main_dev8_inR32[106:7], zll_main_dev8_inR32[6:0], zll_main_dev8_outR32);
  assign zll_main_dev8_inR33 = {main_dev1_in[99:0], 7'h21};
  ZLL_Main_dev8  instR333 (zll_main_dev8_inR33[106:7], zll_main_dev8_inR33[6:0], zll_main_dev8_outR33);
  assign zll_main_dev8_inR34 = {main_dev1_in[99:0], 7'h22};
  ZLL_Main_dev8  instR334 (zll_main_dev8_inR34[106:7], zll_main_dev8_inR34[6:0], zll_main_dev8_outR34);
  assign zll_main_dev8_inR35 = {main_dev1_in[99:0], 7'h23};
  ZLL_Main_dev8  instR335 (zll_main_dev8_inR35[106:7], zll_main_dev8_inR35[6:0], zll_main_dev8_outR35);
  assign zll_main_dev8_inR36 = {main_dev1_in[99:0], 7'h24};
  ZLL_Main_dev8  instR336 (zll_main_dev8_inR36[106:7], zll_main_dev8_inR36[6:0], zll_main_dev8_outR36);
  assign zll_main_dev8_inR37 = {main_dev1_in[99:0], 7'h25};
  ZLL_Main_dev8  instR337 (zll_main_dev8_inR37[106:7], zll_main_dev8_inR37[6:0], zll_main_dev8_outR37);
  assign zll_main_dev8_inR38 = {main_dev1_in[99:0], 7'h26};
  ZLL_Main_dev8  instR338 (zll_main_dev8_inR38[106:7], zll_main_dev8_inR38[6:0], zll_main_dev8_outR38);
  assign zll_main_dev8_inR39 = {main_dev1_in[99:0], 7'h27};
  ZLL_Main_dev8  instR339 (zll_main_dev8_inR39[106:7], zll_main_dev8_inR39[6:0], zll_main_dev8_outR39);
  assign zll_main_dev8_inR40 = {main_dev1_in[99:0], 7'h28};
  ZLL_Main_dev8  instR340 (zll_main_dev8_inR40[106:7], zll_main_dev8_inR40[6:0], zll_main_dev8_outR40);
  assign zll_main_dev8_inR41 = {main_dev1_in[99:0], 7'h29};
  ZLL_Main_dev8  instR341 (zll_main_dev8_inR41[106:7], zll_main_dev8_inR41[6:0], zll_main_dev8_outR41);
  assign zll_main_dev8_inR42 = {main_dev1_in[99:0], 7'h2a};
  ZLL_Main_dev8  instR342 (zll_main_dev8_inR42[106:7], zll_main_dev8_inR42[6:0], zll_main_dev8_outR42);
  assign zll_main_dev8_inR43 = {main_dev1_in[99:0], 7'h2b};
  ZLL_Main_dev8  instR343 (zll_main_dev8_inR43[106:7], zll_main_dev8_inR43[6:0], zll_main_dev8_outR43);
  assign zll_main_dev8_inR44 = {main_dev1_in[99:0], 7'h2c};
  ZLL_Main_dev8  instR344 (zll_main_dev8_inR44[106:7], zll_main_dev8_inR44[6:0], zll_main_dev8_outR44);
  assign zll_main_dev8_inR45 = {main_dev1_in[99:0], 7'h2d};
  ZLL_Main_dev8  instR345 (zll_main_dev8_inR45[106:7], zll_main_dev8_inR45[6:0], zll_main_dev8_outR45);
  assign zll_main_dev8_inR46 = {main_dev1_in[99:0], 7'h2e};
  ZLL_Main_dev8  instR346 (zll_main_dev8_inR46[106:7], zll_main_dev8_inR46[6:0], zll_main_dev8_outR46);
  assign zll_main_dev8_inR47 = {main_dev1_in[99:0], 7'h2f};
  ZLL_Main_dev8  instR347 (zll_main_dev8_inR47[106:7], zll_main_dev8_inR47[6:0], zll_main_dev8_outR47);
  assign zll_main_dev8_inR48 = {main_dev1_in[99:0], 7'h30};
  ZLL_Main_dev8  instR348 (zll_main_dev8_inR48[106:7], zll_main_dev8_inR48[6:0], zll_main_dev8_outR48);
  assign zll_main_dev8_inR49 = {main_dev1_in[99:0], 7'h31};
  ZLL_Main_dev8  instR349 (zll_main_dev8_inR49[106:7], zll_main_dev8_inR49[6:0], zll_main_dev8_outR49);
  assign zll_main_dev8_inR50 = {main_dev1_in[99:0], 7'h32};
  ZLL_Main_dev8  instR350 (zll_main_dev8_inR50[106:7], zll_main_dev8_inR50[6:0], zll_main_dev8_outR50);
  assign zll_main_dev8_inR51 = {main_dev1_in[99:0], 7'h33};
  ZLL_Main_dev8  instR351 (zll_main_dev8_inR51[106:7], zll_main_dev8_inR51[6:0], zll_main_dev8_outR51);
  assign zll_main_dev8_inR52 = {main_dev1_in[99:0], 7'h34};
  ZLL_Main_dev8  instR352 (zll_main_dev8_inR52[106:7], zll_main_dev8_inR52[6:0], zll_main_dev8_outR52);
  assign zll_main_dev8_inR53 = {main_dev1_in[99:0], 7'h35};
  ZLL_Main_dev8  instR353 (zll_main_dev8_inR53[106:7], zll_main_dev8_inR53[6:0], zll_main_dev8_outR53);
  assign zll_main_dev8_inR54 = {main_dev1_in[99:0], 7'h36};
  ZLL_Main_dev8  instR354 (zll_main_dev8_inR54[106:7], zll_main_dev8_inR54[6:0], zll_main_dev8_outR54);
  assign zll_main_dev8_inR55 = {main_dev1_in[99:0], 7'h37};
  ZLL_Main_dev8  instR355 (zll_main_dev8_inR55[106:7], zll_main_dev8_inR55[6:0], zll_main_dev8_outR55);
  assign zll_main_dev8_inR56 = {main_dev1_in[99:0], 7'h38};
  ZLL_Main_dev8  instR356 (zll_main_dev8_inR56[106:7], zll_main_dev8_inR56[6:0], zll_main_dev8_outR56);
  assign zll_main_dev8_inR57 = {main_dev1_in[99:0], 7'h39};
  ZLL_Main_dev8  instR357 (zll_main_dev8_inR57[106:7], zll_main_dev8_inR57[6:0], zll_main_dev8_outR57);
  assign zll_main_dev8_inR58 = {main_dev1_in[99:0], 7'h3a};
  ZLL_Main_dev8  instR358 (zll_main_dev8_inR58[106:7], zll_main_dev8_inR58[6:0], zll_main_dev8_outR58);
  assign zll_main_dev8_inR59 = {main_dev1_in[99:0], 7'h3b};
  ZLL_Main_dev8  instR359 (zll_main_dev8_inR59[106:7], zll_main_dev8_inR59[6:0], zll_main_dev8_outR59);
  assign zll_main_dev8_inR60 = {main_dev1_in[99:0], 7'h3c};
  ZLL_Main_dev8  instR360 (zll_main_dev8_inR60[106:7], zll_main_dev8_inR60[6:0], zll_main_dev8_outR60);
  assign zll_main_dev8_inR61 = {main_dev1_in[99:0], 7'h3d};
  ZLL_Main_dev8  instR361 (zll_main_dev8_inR61[106:7], zll_main_dev8_inR61[6:0], zll_main_dev8_outR61);
  assign zll_main_dev8_inR62 = {main_dev1_in[99:0], 7'h3e};
  ZLL_Main_dev8  instR362 (zll_main_dev8_inR62[106:7], zll_main_dev8_inR62[6:0], zll_main_dev8_outR62);
  assign zll_main_dev8_inR63 = {main_dev1_in[99:0], 7'h3f};
  ZLL_Main_dev8  instR363 (zll_main_dev8_inR63[106:7], zll_main_dev8_inR63[6:0], zll_main_dev8_outR63);
  assign zll_main_dev8_inR64 = {main_dev1_in[99:0], 7'h40};
  ZLL_Main_dev8  instR364 (zll_main_dev8_inR64[106:7], zll_main_dev8_inR64[6:0], zll_main_dev8_outR64);
  assign zll_main_dev8_inR65 = {main_dev1_in[99:0], 7'h41};
  ZLL_Main_dev8  instR365 (zll_main_dev8_inR65[106:7], zll_main_dev8_inR65[6:0], zll_main_dev8_outR65);
  assign zll_main_dev8_inR66 = {main_dev1_in[99:0], 7'h42};
  ZLL_Main_dev8  instR366 (zll_main_dev8_inR66[106:7], zll_main_dev8_inR66[6:0], zll_main_dev8_outR66);
  assign zll_main_dev8_inR67 = {main_dev1_in[99:0], 7'h43};
  ZLL_Main_dev8  instR367 (zll_main_dev8_inR67[106:7], zll_main_dev8_inR67[6:0], zll_main_dev8_outR67);
  assign zll_main_dev8_inR68 = {main_dev1_in[99:0], 7'h44};
  ZLL_Main_dev8  instR368 (zll_main_dev8_inR68[106:7], zll_main_dev8_inR68[6:0], zll_main_dev8_outR68);
  assign zll_main_dev8_inR69 = {main_dev1_in[99:0], 7'h45};
  ZLL_Main_dev8  instR369 (zll_main_dev8_inR69[106:7], zll_main_dev8_inR69[6:0], zll_main_dev8_outR69);
  assign zll_main_dev8_inR70 = {main_dev1_in[99:0], 7'h46};
  ZLL_Main_dev8  instR370 (zll_main_dev8_inR70[106:7], zll_main_dev8_inR70[6:0], zll_main_dev8_outR70);
  assign zll_main_dev8_inR71 = {main_dev1_in[99:0], 7'h47};
  ZLL_Main_dev8  instR371 (zll_main_dev8_inR71[106:7], zll_main_dev8_inR71[6:0], zll_main_dev8_outR71);
  assign zll_main_dev8_inR72 = {main_dev1_in[99:0], 7'h48};
  ZLL_Main_dev8  instR372 (zll_main_dev8_inR72[106:7], zll_main_dev8_inR72[6:0], zll_main_dev8_outR72);
  assign zll_main_dev8_inR73 = {main_dev1_in[99:0], 7'h49};
  ZLL_Main_dev8  instR373 (zll_main_dev8_inR73[106:7], zll_main_dev8_inR73[6:0], zll_main_dev8_outR73);
  assign zll_main_dev8_inR74 = {main_dev1_in[99:0], 7'h4a};
  ZLL_Main_dev8  instR374 (zll_main_dev8_inR74[106:7], zll_main_dev8_inR74[6:0], zll_main_dev8_outR74);
  assign zll_main_dev8_inR75 = {main_dev1_in[99:0], 7'h4b};
  ZLL_Main_dev8  instR375 (zll_main_dev8_inR75[106:7], zll_main_dev8_inR75[6:0], zll_main_dev8_outR75);
  assign zll_main_dev8_inR76 = {main_dev1_in[99:0], 7'h4c};
  ZLL_Main_dev8  instR376 (zll_main_dev8_inR76[106:7], zll_main_dev8_inR76[6:0], zll_main_dev8_outR76);
  assign zll_main_dev8_inR77 = {main_dev1_in[99:0], 7'h4d};
  ZLL_Main_dev8  instR377 (zll_main_dev8_inR77[106:7], zll_main_dev8_inR77[6:0], zll_main_dev8_outR77);
  assign zll_main_dev8_inR78 = {main_dev1_in[99:0], 7'h4e};
  ZLL_Main_dev8  instR378 (zll_main_dev8_inR78[106:7], zll_main_dev8_inR78[6:0], zll_main_dev8_outR78);
  assign zll_main_dev8_inR79 = {main_dev1_in[99:0], 7'h4f};
  ZLL_Main_dev8  instR379 (zll_main_dev8_inR79[106:7], zll_main_dev8_inR79[6:0], zll_main_dev8_outR79);
  assign zll_main_dev8_inR80 = {main_dev1_in[99:0], 7'h50};
  ZLL_Main_dev8  instR380 (zll_main_dev8_inR80[106:7], zll_main_dev8_inR80[6:0], zll_main_dev8_outR80);
  assign zll_main_dev8_inR81 = {main_dev1_in[99:0], 7'h51};
  ZLL_Main_dev8  instR381 (zll_main_dev8_inR81[106:7], zll_main_dev8_inR81[6:0], zll_main_dev8_outR81);
  assign zll_main_dev8_inR82 = {main_dev1_in[99:0], 7'h52};
  ZLL_Main_dev8  instR382 (zll_main_dev8_inR82[106:7], zll_main_dev8_inR82[6:0], zll_main_dev8_outR82);
  assign zll_main_dev8_inR83 = {main_dev1_in[99:0], 7'h53};
  ZLL_Main_dev8  instR383 (zll_main_dev8_inR83[106:7], zll_main_dev8_inR83[6:0], zll_main_dev8_outR83);
  assign zll_main_dev8_inR84 = {main_dev1_in[99:0], 7'h54};
  ZLL_Main_dev8  instR384 (zll_main_dev8_inR84[106:7], zll_main_dev8_inR84[6:0], zll_main_dev8_outR84);
  assign zll_main_dev8_inR85 = {main_dev1_in[99:0], 7'h55};
  ZLL_Main_dev8  instR385 (zll_main_dev8_inR85[106:7], zll_main_dev8_inR85[6:0], zll_main_dev8_outR85);
  assign zll_main_dev8_inR86 = {main_dev1_in[99:0], 7'h56};
  ZLL_Main_dev8  instR386 (zll_main_dev8_inR86[106:7], zll_main_dev8_inR86[6:0], zll_main_dev8_outR86);
  assign zll_main_dev8_inR87 = {main_dev1_in[99:0], 7'h57};
  ZLL_Main_dev8  instR387 (zll_main_dev8_inR87[106:7], zll_main_dev8_inR87[6:0], zll_main_dev8_outR87);
  assign zll_main_dev8_inR88 = {main_dev1_in[99:0], 7'h58};
  ZLL_Main_dev8  instR388 (zll_main_dev8_inR88[106:7], zll_main_dev8_inR88[6:0], zll_main_dev8_outR88);
  assign zll_main_dev8_inR89 = {main_dev1_in[99:0], 7'h59};
  ZLL_Main_dev8  instR389 (zll_main_dev8_inR89[106:7], zll_main_dev8_inR89[6:0], zll_main_dev8_outR89);
  assign zll_main_dev8_inR90 = {main_dev1_in[99:0], 7'h5a};
  ZLL_Main_dev8  instR390 (zll_main_dev8_inR90[106:7], zll_main_dev8_inR90[6:0], zll_main_dev8_outR90);
  assign zll_main_dev8_inR91 = {main_dev1_in[99:0], 7'h5b};
  ZLL_Main_dev8  instR391 (zll_main_dev8_inR91[106:7], zll_main_dev8_inR91[6:0], zll_main_dev8_outR91);
  assign zll_main_dev8_inR92 = {main_dev1_in[99:0], 7'h5c};
  ZLL_Main_dev8  instR392 (zll_main_dev8_inR92[106:7], zll_main_dev8_inR92[6:0], zll_main_dev8_outR92);
  assign zll_main_dev8_inR93 = {main_dev1_in[99:0], 7'h5d};
  ZLL_Main_dev8  instR393 (zll_main_dev8_inR93[106:7], zll_main_dev8_inR93[6:0], zll_main_dev8_outR93);
  assign zll_main_dev8_inR94 = {main_dev1_in[99:0], 7'h5e};
  ZLL_Main_dev8  instR394 (zll_main_dev8_inR94[106:7], zll_main_dev8_inR94[6:0], zll_main_dev8_outR94);
  assign zll_main_dev8_inR95 = {main_dev1_in[99:0], 7'h5f};
  ZLL_Main_dev8  instR395 (zll_main_dev8_inR95[106:7], zll_main_dev8_inR95[6:0], zll_main_dev8_outR95);
  assign zll_main_dev8_inR96 = {main_dev1_in[99:0], 7'h60};
  ZLL_Main_dev8  instR396 (zll_main_dev8_inR96[106:7], zll_main_dev8_inR96[6:0], zll_main_dev8_outR96);
  assign zll_main_dev8_inR97 = {main_dev1_in[99:0], 7'h61};
  ZLL_Main_dev8  instR397 (zll_main_dev8_inR97[106:7], zll_main_dev8_inR97[6:0], zll_main_dev8_outR97);
  assign zll_main_dev8_inR98 = {main_dev1_in[99:0], 7'h62};
  ZLL_Main_dev8  instR398 (zll_main_dev8_inR98[106:7], zll_main_dev8_inR98[6:0], zll_main_dev8_outR98);
  assign zll_main_dev8_inR99 = {main_dev1_in[99:0], 7'h63};
  ZLL_Main_dev8  instR399 (zll_main_dev8_inR99[106:7], zll_main_dev8_inR99[6:0], zll_main_dev8_outR99);
  assign {__continue, __out0, __out1, __out2, __out3, __resumption_tag_next} = {zll_main_dev20_out, zll_main_dev20_outR1, zll_main_dev20_outR2, zll_main_dev20_outR3, zll_main_dev20_outR4, zll_main_dev20_outR5, zll_main_dev20_outR6, zll_main_dev20_outR7, zll_main_dev20_outR8, zll_main_dev20_outR9, zll_main_dev20_outR10, zll_main_dev20_outR11, zll_main_dev20_outR12, zll_main_dev20_outR13, zll_main_dev20_outR14, zll_main_dev20_outR15, zll_main_dev20_outR16, zll_main_dev20_outR17, zll_main_dev20_outR18, zll_main_dev20_outR19, zll_main_dev20_outR20, zll_main_dev20_outR21, zll_main_dev20_outR22, zll_main_dev20_outR23, zll_main_dev20_outR24, zll_main_dev20_outR25, zll_main_dev20_outR26, zll_main_dev20_outR27, zll_main_dev20_outR28, zll_main_dev20_outR29, zll_main_dev20_outR30, zll_main_dev20_outR31, zll_main_dev20_outR32, zll_main_dev20_outR33, zll_main_dev20_outR34, zll_main_dev20_outR35, zll_main_dev20_outR36, zll_main_dev20_outR37, zll_main_dev20_outR38, zll_main_dev20_outR39, zll_main_dev20_outR40, zll_main_dev20_outR41, zll_main_dev20_outR42, zll_main_dev20_outR43, zll_main_dev20_outR44, zll_main_dev20_outR45, zll_main_dev20_outR46, zll_main_dev20_outR47, zll_main_dev20_outR48, zll_main_dev20_outR49, zll_main_dev20_outR50, zll_main_dev20_outR51, zll_main_dev20_outR52, zll_main_dev20_outR53, zll_main_dev20_outR54, zll_main_dev20_outR55, zll_main_dev20_outR56, zll_main_dev20_outR57, zll_main_dev20_outR58, zll_main_dev20_outR59, zll_main_dev20_outR60, zll_main_dev20_outR61, zll_main_dev20_outR62, zll_main_dev20_outR63, zll_main_dev20_outR64, zll_main_dev20_outR65, zll_main_dev20_outR66, zll_main_dev20_outR67, zll_main_dev20_outR68, zll_main_dev20_outR69, zll_main_dev20_outR70, zll_main_dev20_outR71, zll_main_dev20_outR72, zll_main_dev20_outR73, zll_main_dev20_outR74, zll_main_dev20_outR75, zll_main_dev20_outR76, zll_main_dev20_outR77, zll_main_dev20_outR78, zll_main_dev20_outR79, zll_main_dev20_outR80, zll_main_dev20_outR81, zll_main_dev20_outR82, zll_main_dev20_outR83, zll_main_dev20_outR84, zll_main_dev20_outR85, zll_main_dev20_outR86, zll_main_dev20_outR87, zll_main_dev20_outR88, zll_main_dev20_outR89, zll_main_dev20_outR90, zll_main_dev20_outR91, zll_main_dev20_outR92, zll_main_dev20_outR93, zll_main_dev20_outR94, zll_main_dev20_outR95, zll_main_dev20_outR96, zll_main_dev20_outR97, zll_main_dev20_outR98, zll_main_dev20_outR99, zll_main_dev12_out, zll_main_dev12_outR1, zll_main_dev12_outR2, zll_main_dev12_outR3, zll_main_dev12_outR4, zll_main_dev12_outR5, zll_main_dev12_outR6, zll_main_dev12_outR7, zll_main_dev12_outR8, zll_main_dev12_outR9, zll_main_dev12_outR10, zll_main_dev12_outR11, zll_main_dev12_outR12, zll_main_dev12_outR13, zll_main_dev12_outR14, zll_main_dev12_outR15, zll_main_dev12_outR16, zll_main_dev12_outR17, zll_main_dev12_outR18, zll_main_dev12_outR19, zll_main_dev12_outR20, zll_main_dev12_outR21, zll_main_dev12_outR22, zll_main_dev12_outR23, zll_main_dev12_outR24, zll_main_dev12_outR25, zll_main_dev12_outR26, zll_main_dev12_outR27, zll_main_dev12_outR28, zll_main_dev12_outR29, zll_main_dev12_outR30, zll_main_dev12_outR31, zll_main_dev12_outR32, zll_main_dev12_outR33, zll_main_dev12_outR34, zll_main_dev12_outR35, zll_main_dev12_outR36, zll_main_dev12_outR37, zll_main_dev12_outR38, zll_main_dev12_outR39, zll_main_dev12_outR40, zll_main_dev12_outR41, zll_main_dev12_outR42, zll_main_dev12_outR43, zll_main_dev12_outR44, zll_main_dev12_outR45, zll_main_dev12_outR46, zll_main_dev12_outR47, zll_main_dev12_outR48, zll_main_dev12_outR49, zll_main_dev12_outR50, zll_main_dev12_outR51, zll_main_dev12_outR52, zll_main_dev12_outR53, zll_main_dev12_outR54, zll_main_dev12_outR55, zll_main_dev12_outR56, zll_main_dev12_outR57, zll_main_dev12_outR58, zll_main_dev12_outR59, zll_main_dev12_outR60, zll_main_dev12_outR61, zll_main_dev12_outR62, zll_main_dev12_outR63, zll_main_dev12_outR64, zll_main_dev12_outR65, zll_main_dev12_outR66, zll_main_dev12_outR67, zll_main_dev12_outR68, zll_main_dev12_outR69, zll_main_dev12_outR70, zll_main_dev12_outR71, zll_main_dev12_outR72, zll_main_dev12_outR73, zll_main_dev12_outR74, zll_main_dev12_outR75, zll_main_dev12_outR76, zll_main_dev12_outR77, zll_main_dev12_outR78, zll_main_dev12_outR79, zll_main_dev12_outR80, zll_main_dev12_outR81, zll_main_dev12_outR82, zll_main_dev12_outR83, zll_main_dev12_outR84, zll_main_dev12_outR85, zll_main_dev12_outR86, zll_main_dev12_outR87, zll_main_dev12_outR88, zll_main_dev12_outR89, zll_main_dev12_outR90, zll_main_dev12_outR91, zll_main_dev12_outR92, zll_main_dev12_outR93, zll_main_dev12_outR94, zll_main_dev12_outR95, zll_main_dev12_outR96, zll_main_dev12_outR97, zll_main_dev12_outR98, zll_main_dev12_outR99, zll_main_dev15_out, zll_main_dev15_outR1, zll_main_dev15_outR2, zll_main_dev15_outR3, zll_main_dev15_outR4, zll_main_dev15_outR5, zll_main_dev15_outR6, zll_main_dev15_outR7, zll_main_dev15_outR8, zll_main_dev15_outR9, zll_main_dev15_outR10, zll_main_dev15_outR11, zll_main_dev15_outR12, zll_main_dev15_outR13, zll_main_dev15_outR14, zll_main_dev15_outR15, zll_main_dev15_outR16, zll_main_dev15_outR17, zll_main_dev15_outR18, zll_main_dev15_outR19, zll_main_dev15_outR20, zll_main_dev15_outR21, zll_main_dev15_outR22, zll_main_dev15_outR23, zll_main_dev15_outR24, zll_main_dev15_outR25, zll_main_dev15_outR26, zll_main_dev15_outR27, zll_main_dev15_outR28, zll_main_dev15_outR29, zll_main_dev15_outR30, zll_main_dev15_outR31, zll_main_dev15_outR32, zll_main_dev15_outR33, zll_main_dev15_outR34, zll_main_dev15_outR35, zll_main_dev15_outR36, zll_main_dev15_outR37, zll_main_dev15_outR38, zll_main_dev15_outR39, zll_main_dev15_outR40, zll_main_dev15_outR41, zll_main_dev15_outR42, zll_main_dev15_outR43, zll_main_dev15_outR44, zll_main_dev15_outR45, zll_main_dev15_outR46, zll_main_dev15_outR47, zll_main_dev15_outR48, zll_main_dev15_outR49, zll_main_dev15_outR50, zll_main_dev15_outR51, zll_main_dev15_outR52, zll_main_dev15_outR53, zll_main_dev15_outR54, zll_main_dev15_outR55, zll_main_dev15_outR56, zll_main_dev15_outR57, zll_main_dev15_outR58, zll_main_dev15_outR59, zll_main_dev15_outR60, zll_main_dev15_outR61, zll_main_dev15_outR62, zll_main_dev15_outR63, zll_main_dev15_outR64, zll_main_dev15_outR65, zll_main_dev15_outR66, zll_main_dev15_outR67, zll_main_dev15_outR68, zll_main_dev15_outR69, zll_main_dev15_outR70, zll_main_dev15_outR71, zll_main_dev15_outR72, zll_main_dev15_outR73, zll_main_dev15_outR74, zll_main_dev15_outR75, zll_main_dev15_outR76, zll_main_dev15_outR77, zll_main_dev15_outR78, zll_main_dev15_outR79, zll_main_dev15_outR80, zll_main_dev15_outR81, zll_main_dev15_outR82, zll_main_dev15_outR83, zll_main_dev15_outR84, zll_main_dev15_outR85, zll_main_dev15_outR86, zll_main_dev15_outR87, zll_main_dev15_outR88, zll_main_dev15_outR89, zll_main_dev15_outR90, zll_main_dev15_outR91, zll_main_dev15_outR92, zll_main_dev15_outR93, zll_main_dev15_outR94, zll_main_dev15_outR95, zll_main_dev15_outR96, zll_main_dev15_outR97, zll_main_dev15_outR98, zll_main_dev15_outR99, zll_main_dev8_out, zll_main_dev8_outR1, zll_main_dev8_outR2, zll_main_dev8_outR3, zll_main_dev8_outR4, zll_main_dev8_outR5, zll_main_dev8_outR6, zll_main_dev8_outR7, zll_main_dev8_outR8, zll_main_dev8_outR9, zll_main_dev8_outR10, zll_main_dev8_outR11, zll_main_dev8_outR12, zll_main_dev8_outR13, zll_main_dev8_outR14, zll_main_dev8_outR15, zll_main_dev8_outR16, zll_main_dev8_outR17, zll_main_dev8_outR18, zll_main_dev8_outR19, zll_main_dev8_outR20, zll_main_dev8_outR21, zll_main_dev8_outR22, zll_main_dev8_outR23, zll_main_dev8_outR24, zll_main_dev8_outR25, zll_main_dev8_outR26, zll_main_dev8_outR27, zll_main_dev8_outR28, zll_main_dev8_outR29, zll_main_dev8_outR30, zll_main_dev8_outR31, zll_main_dev8_outR32, zll_main_dev8_outR33, zll_main_dev8_outR34, zll_main_dev8_outR35, zll_main_dev8_outR36, zll_main_dev8_outR37, zll_main_dev8_outR38, zll_main_dev8_outR39, zll_main_dev8_outR40, zll_main_dev8_outR41, zll_main_dev8_outR42, zll_main_dev8_outR43, zll_main_dev8_outR44, zll_main_dev8_outR45, zll_main_dev8_outR46, zll_main_dev8_outR47, zll_main_dev8_outR48, zll_main_dev8_outR49, zll_main_dev8_outR50, zll_main_dev8_outR51, zll_main_dev8_outR52, zll_main_dev8_outR53, zll_main_dev8_outR54, zll_main_dev8_outR55, zll_main_dev8_outR56, zll_main_dev8_outR57, zll_main_dev8_outR58, zll_main_dev8_outR59, zll_main_dev8_outR60, zll_main_dev8_outR61, zll_main_dev8_outR62, zll_main_dev8_outR63, zll_main_dev8_outR64, zll_main_dev8_outR65, zll_main_dev8_outR66, zll_main_dev8_outR67, zll_main_dev8_outR68, zll_main_dev8_outR69, zll_main_dev8_outR70, zll_main_dev8_outR71, zll_main_dev8_outR72, zll_main_dev8_outR73, zll_main_dev8_outR74, zll_main_dev8_outR75, zll_main_dev8_outR76, zll_main_dev8_outR77, zll_main_dev8_outR78, zll_main_dev8_outR79, zll_main_dev8_outR80, zll_main_dev8_outR81, zll_main_dev8_outR82, zll_main_dev8_outR83, zll_main_dev8_outR84, zll_main_dev8_outR85, zll_main_dev8_outR86, zll_main_dev8_outR87, zll_main_dev8_outR88, zll_main_dev8_outR89, zll_main_dev8_outR90, zll_main_dev8_outR91, zll_main_dev8_outR92, zll_main_dev8_outR93, zll_main_dev8_outR94, zll_main_dev8_outR95, zll_main_dev8_outR96, zll_main_dev8_outR97, zll_main_dev8_outR98, zll_main_dev8_outR99};
  initial __resumption_tag <= {7'h64{1'h0}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      __resumption_tag <= {7'h64{1'h0}};
    end else begin
      __resumption_tag <= __resumption_tag_next;
    end
  end
endmodule

module ZLL_Main_dev20 (input logic [99:0] arg0,
  input logic [6:0] arg1,
  output logic [0:0] res);
  logic [6:0] resize_in;
  logic [127:0] resize_inR1;
  logic [0:0] msbit_in;
  logic [0:0] rewire_prelude_not_in;
  logic [0:0] rewire_prelude_not_out;
  logic [6:0] resize_inR2;
  logic [127:0] resize_inR3;
  logic [0:0] msbit_inR1;
  logic [0:0] rewire_prelude_not_inR1;
  logic [0:0] rewire_prelude_not_outR1;
  logic [107:0] zll_main_dev4_in;
  logic [99:0] main_x2_in;
  logic [99:0] main_x2_out;
  logic [99:0] resize_inR4;
  logic [6:0] resize_inR5;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR6;
  logic [6:0] resize_inR7;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR8;
  logic [6:0] resize_inR9;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR10;
  logic [107:0] zll_main_dev11_in;
  logic [99:0] resize_inR11;
  logic [6:0] resize_inR12;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR13;
  logic [6:0] resize_inR14;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [127:0] resize_inR15;
  assign resize_in = arg1;
  assign resize_inR1 = 128'(resize_in[6:0]);
  assign msbit_in = resize_inR1[0];
  assign rewire_prelude_not_in = msbit_in[0];
  ReWire_Prelude_not  inst (rewire_prelude_not_in[0], rewire_prelude_not_out);
  assign resize_inR2 = arg1;
  assign resize_inR3 = 128'(resize_inR2[6:0]);
  assign msbit_inR1 = resize_inR3[0];
  assign rewire_prelude_not_inR1 = msbit_inR1[0];
  ReWire_Prelude_not  instR1 (rewire_prelude_not_inR1[0], rewire_prelude_not_outR1);
  assign zll_main_dev4_in = {arg0, arg1, rewire_prelude_not_outR1};
  assign main_x2_in = zll_main_dev4_in[107:8];
  Main_x2  instR2 (main_x2_in[99:0], main_x2_out);
  assign resize_inR4 = main_x2_out;
  assign resize_inR5 = zll_main_dev4_in[7:1];
  assign binop_in = {128'(resize_inR5[6:0]), 128'h1};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h64};
  assign resize_inR6 = binop_inR1[255:128] % binop_inR1[127:0];
  assign resize_inR7 = resize_inR6[6:0];
  assign binop_inR2 = {128'(resize_inR7[6:0]), 128'h2};
  assign binop_inR3 = {binop_inR2[255:128] / binop_inR2[127:0], 128'h64};
  assign resize_inR8 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR9 = resize_inR8[6:0];
  assign binop_inR4 = {128'h64, 128'(resize_inR9[6:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h1};
  assign binop_inR7 = {128'(resize_inR4[99:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR10 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign zll_main_dev11_in = {arg0, arg1, rewire_prelude_not_out};
  assign resize_inR11 = zll_main_dev11_in[107:8];
  assign resize_inR12 = zll_main_dev11_in[7:1];
  assign binop_inR8 = {128'(resize_inR12[6:0]), 128'h2};
  assign binop_inR9 = {binop_inR8[255:128] / binop_inR8[127:0], 128'h64};
  assign resize_inR13 = binop_inR9[255:128] % binop_inR9[127:0];
  assign resize_inR14 = resize_inR13[6:0];
  assign binop_inR10 = {128'h64, 128'(resize_inR14[6:0])};
  assign binop_inR11 = {binop_inR10[255:128] - binop_inR10[127:0], 128'h1};
  assign binop_inR12 = {binop_inR11[255:128] - binop_inR11[127:0], 128'h1};
  assign binop_inR13 = {128'(resize_inR11[99:0]), binop_inR12[255:128] * binop_inR12[127:0]};
  assign resize_inR15 = binop_inR13[255:128] >> binop_inR13[127:0];
  assign res = (zll_main_dev11_in[0] == 1'h1) ? resize_inR15[0] : resize_inR10[0];
endmodule

module ReWire_Prelude_not (input logic [0:0] arg0,
  output logic [0:0] res);
  logic [0:0] lit_in;
  assign lit_in = arg0;
  assign res = (lit_in[0] == 1'h1) ? 1'h0 : 1'h1;
endmodule

module ZLL_Main_dev15 (input logic [99:0] arg0,
  input logic [6:0] arg1,
  output logic [0:0] res);
  logic [6:0] resize_in;
  logic [255:0] binop_in;
  logic [6:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [107:0] zll_main_dev10_in;
  logic [99:0] main_x2_in;
  logic [99:0] main_x2_out;
  logic [99:0] resize_inR2;
  logic [6:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [6:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [6:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR8;
  logic [107:0] zll_main_dev14_in;
  logic [99:0] resize_inR9;
  logic [6:0] resize_inR10;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR11;
  logic [6:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR13;
  assign resize_in = arg1;
  assign binop_in = {128'(resize_in[6:0]), 128'h31};
  assign resize_inR1 = arg1;
  assign binop_inR1 = {128'(resize_inR1[6:0]), 128'h31};
  assign zll_main_dev10_in = {arg0, arg1, binop_inR1[255:128] < binop_inR1[127:0]};
  assign main_x2_in = zll_main_dev10_in[107:8];
  Main_x2  inst (main_x2_in[99:0], main_x2_out);
  assign resize_inR2 = main_x2_out;
  assign resize_inR3 = zll_main_dev10_in[7:1];
  assign binop_inR2 = {128'(resize_inR3[6:0]), 128'h31};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h64};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[6:0];
  assign binop_inR4 = {128'(resize_inR5[6:0]), 128'h2};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h64};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[6:0];
  assign binop_inR6 = {128'h64, 128'(resize_inR7[6:0])};
  assign binop_inR7 = {binop_inR6[255:128] - binop_inR6[127:0], 128'h1};
  assign binop_inR8 = {binop_inR7[255:128] - binop_inR7[127:0], 128'h1};
  assign binop_inR9 = {128'(resize_inR2[99:0]), binop_inR8[255:128] * binop_inR8[127:0]};
  assign resize_inR8 = binop_inR9[255:128] >> binop_inR9[127:0];
  assign zll_main_dev14_in = {arg0, arg1, binop_in[255:128] < binop_in[127:0]};
  assign resize_inR9 = zll_main_dev14_in[107:8];
  assign resize_inR10 = zll_main_dev14_in[7:1];
  assign binop_inR10 = {128'(resize_inR10[6:0]), 128'h2};
  assign binop_inR11 = {binop_inR10[255:128] * binop_inR10[127:0], 128'h64};
  assign resize_inR11 = binop_inR11[255:128] % binop_inR11[127:0];
  assign resize_inR12 = resize_inR11[6:0];
  assign binop_inR12 = {128'h64, 128'(resize_inR12[6:0])};
  assign binop_inR13 = {binop_inR12[255:128] - binop_inR12[127:0], 128'h1};
  assign binop_inR14 = {binop_inR13[255:128] - binop_inR13[127:0], 128'h1};
  assign binop_inR15 = {128'(resize_inR9[99:0]), binop_inR14[255:128] * binop_inR14[127:0]};
  assign resize_inR13 = binop_inR15[255:128] >> binop_inR15[127:0];
  assign res = (zll_main_dev14_in[0] == 1'h1) ? resize_inR13[0] : resize_inR8[0];
endmodule

module ZLL_Main_dev12 (input logic [99:0] arg0,
  input logic [6:0] arg1,
  output logic [0:0] res);
  logic [6:0] resize_in;
  logic [127:0] resize_inR1;
  logic [0:0] msbit_in;
  logic [0:0] rewire_prelude_not_in;
  logic [0:0] rewire_prelude_not_out;
  logic [6:0] resize_inR2;
  logic [127:0] resize_inR3;
  logic [0:0] msbit_inR1;
  logic [0:0] rewire_prelude_not_inR1;
  logic [0:0] rewire_prelude_not_outR1;
  logic [107:0] zll_main_dev13_in;
  logic [99:0] main_x2_in;
  logic [99:0] main_x2_out;
  logic [99:0] resize_inR4;
  logic [6:0] resize_inR5;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR6;
  logic [6:0] resize_inR7;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR8;
  logic [6:0] resize_inR9;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR10;
  logic [6:0] resize_inR11;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR12;
  logic [107:0] zll_main_dev18_in;
  logic [99:0] resize_inR13;
  logic [6:0] resize_inR14;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR15;
  logic [6:0] resize_inR16;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [127:0] resize_inR17;
  logic [6:0] resize_inR18;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [255:0] binop_inR16;
  logic [255:0] binop_inR17;
  logic [127:0] resize_inR19;
  assign resize_in = arg1;
  assign resize_inR1 = 128'(resize_in[6:0]);
  assign msbit_in = resize_inR1[0];
  assign rewire_prelude_not_in = msbit_in[0];
  ReWire_Prelude_not  inst (rewire_prelude_not_in[0], rewire_prelude_not_out);
  assign resize_inR2 = arg1;
  assign resize_inR3 = 128'(resize_inR2[6:0]);
  assign msbit_inR1 = resize_inR3[0];
  assign rewire_prelude_not_inR1 = msbit_inR1[0];
  ReWire_Prelude_not  instR1 (rewire_prelude_not_inR1[0], rewire_prelude_not_outR1);
  assign zll_main_dev13_in = {arg0, arg1, rewire_prelude_not_outR1};
  assign main_x2_in = zll_main_dev13_in[107:8];
  Main_x2  instR2 (main_x2_in[99:0], main_x2_out);
  assign resize_inR4 = main_x2_out;
  assign resize_inR5 = zll_main_dev13_in[7:1];
  assign binop_in = {128'(resize_inR5[6:0]), 128'h1};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h64};
  assign resize_inR6 = binop_inR1[255:128] % binop_inR1[127:0];
  assign resize_inR7 = resize_inR6[6:0];
  assign binop_inR2 = {128'h31, 128'(resize_inR7[6:0])};
  assign binop_inR3 = {binop_inR2[255:128] + binop_inR2[127:0], 128'h64};
  assign resize_inR8 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR9 = resize_inR8[6:0];
  assign binop_inR4 = {128'(resize_inR9[6:0]), 128'h2};
  assign binop_inR5 = {binop_inR4[255:128] / binop_inR4[127:0], 128'h64};
  assign resize_inR10 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR11 = resize_inR10[6:0];
  assign binop_inR6 = {128'h64, 128'(resize_inR11[6:0])};
  assign binop_inR7 = {binop_inR6[255:128] - binop_inR6[127:0], 128'h1};
  assign binop_inR8 = {binop_inR7[255:128] - binop_inR7[127:0], 128'h1};
  assign binop_inR9 = {128'(resize_inR4[99:0]), binop_inR8[255:128] * binop_inR8[127:0]};
  assign resize_inR12 = binop_inR9[255:128] >> binop_inR9[127:0];
  assign zll_main_dev18_in = {arg0, arg1, rewire_prelude_not_out};
  assign resize_inR13 = zll_main_dev18_in[107:8];
  assign resize_inR14 = zll_main_dev18_in[7:1];
  assign binop_inR10 = {128'h31, 128'(resize_inR14[6:0])};
  assign binop_inR11 = {binop_inR10[255:128] + binop_inR10[127:0], 128'h64};
  assign resize_inR15 = binop_inR11[255:128] % binop_inR11[127:0];
  assign resize_inR16 = resize_inR15[6:0];
  assign binop_inR12 = {128'(resize_inR16[6:0]), 128'h2};
  assign binop_inR13 = {binop_inR12[255:128] / binop_inR12[127:0], 128'h64};
  assign resize_inR17 = binop_inR13[255:128] % binop_inR13[127:0];
  assign resize_inR18 = resize_inR17[6:0];
  assign binop_inR14 = {128'h64, 128'(resize_inR18[6:0])};
  assign binop_inR15 = {binop_inR14[255:128] - binop_inR14[127:0], 128'h1};
  assign binop_inR16 = {binop_inR15[255:128] - binop_inR15[127:0], 128'h1};
  assign binop_inR17 = {128'(resize_inR13[99:0]), binop_inR16[255:128] * binop_inR16[127:0]};
  assign resize_inR19 = binop_inR17[255:128] >> binop_inR17[127:0];
  assign res = (zll_main_dev18_in[0] == 1'h1) ? resize_inR19[0] : resize_inR12[0];
endmodule

module ZLL_Main_dev8 (input logic [99:0] arg0,
  input logic [6:0] arg1,
  output logic [0:0] res);
  logic [6:0] resize_in;
  logic [255:0] binop_in;
  logic [6:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [107:0] zll_main_dev21_in;
  logic [99:0] main_x2_in;
  logic [99:0] main_x2_out;
  logic [99:0] resize_inR2;
  logic [6:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [6:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [6:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR8;
  logic [6:0] resize_inR9;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR10;
  logic [107:0] zll_main_dev23_in;
  logic [99:0] resize_inR11;
  logic [6:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [127:0] resize_inR13;
  logic [6:0] resize_inR14;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR15;
  logic [6:0] resize_inR16;
  logic [255:0] binop_inR16;
  logic [255:0] binop_inR17;
  logic [255:0] binop_inR18;
  logic [255:0] binop_inR19;
  logic [127:0] resize_inR17;
  assign resize_in = arg1;
  assign binop_in = {128'(resize_in[6:0]), 128'h31};
  assign resize_inR1 = arg1;
  assign binop_inR1 = {128'(resize_inR1[6:0]), 128'h31};
  assign zll_main_dev21_in = {arg0, arg1, binop_inR1[255:128] < binop_inR1[127:0]};
  assign main_x2_in = zll_main_dev21_in[107:8];
  Main_x2  inst (main_x2_in[99:0], main_x2_out);
  assign resize_inR2 = main_x2_out;
  assign resize_inR3 = zll_main_dev21_in[7:1];
  assign binop_inR2 = {128'(resize_inR3[6:0]), 128'h31};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h64};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[6:0];
  assign binop_inR4 = {128'(resize_inR5[6:0]), 128'h2};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h64};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[6:0];
  assign binop_inR6 = {128'(resize_inR7[6:0]), 128'h1};
  assign binop_inR7 = {binop_inR6[255:128] + binop_inR6[127:0], 128'h64};
  assign resize_inR8 = binop_inR7[255:128] % binop_inR7[127:0];
  assign resize_inR9 = resize_inR8[6:0];
  assign binop_inR8 = {128'h64, 128'(resize_inR9[6:0])};
  assign binop_inR9 = {binop_inR8[255:128] - binop_inR8[127:0], 128'h1};
  assign binop_inR10 = {binop_inR9[255:128] - binop_inR9[127:0], 128'h1};
  assign binop_inR11 = {128'(resize_inR2[99:0]), binop_inR10[255:128] * binop_inR10[127:0]};
  assign resize_inR10 = binop_inR11[255:128] >> binop_inR11[127:0];
  assign zll_main_dev23_in = {arg0, arg1, binop_in[255:128] < binop_in[127:0]};
  assign resize_inR11 = zll_main_dev23_in[107:8];
  assign resize_inR12 = zll_main_dev23_in[7:1];
  assign binop_inR12 = {128'(resize_inR12[6:0]), 128'h2};
  assign binop_inR13 = {binop_inR12[255:128] * binop_inR12[127:0], 128'h64};
  assign resize_inR13 = binop_inR13[255:128] % binop_inR13[127:0];
  assign resize_inR14 = resize_inR13[6:0];
  assign binop_inR14 = {128'(resize_inR14[6:0]), 128'h1};
  assign binop_inR15 = {binop_inR14[255:128] + binop_inR14[127:0], 128'h64};
  assign resize_inR15 = binop_inR15[255:128] % binop_inR15[127:0];
  assign resize_inR16 = resize_inR15[6:0];
  assign binop_inR16 = {128'h64, 128'(resize_inR16[6:0])};
  assign binop_inR17 = {binop_inR16[255:128] - binop_inR16[127:0], 128'h1};
  assign binop_inR18 = {binop_inR17[255:128] - binop_inR17[127:0], 128'h1};
  assign binop_inR19 = {128'(resize_inR11[99:0]), binop_inR18[255:128] * binop_inR18[127:0]};
  assign resize_inR17 = binop_inR19[255:128] >> binop_inR19[127:0];
  assign res = (zll_main_dev23_in[0] == 1'h1) ? resize_inR17[0] : resize_inR10[0];
endmodule

module Main_x2 (input logic [99:0] arg0,
  output logic [99:0] res);
  logic [199:0] binop_in;
  assign binop_in = {arg0, 100'h2};
  assign res = binop_in[199:100] * binop_in[99:0];
endmodule