module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [16:0] __in0,
  output logic [14:0] __out0);
  logic [90:0] zll_pure_dispatch7_in;
  logic [142:0] zll_pure_dispatch7_out;
  logic [90:0] zll_pure_dispatch7_inR1;
  logic [142:0] zll_pure_dispatch7_outR1;
  logic [90:0] zll_pure_dispatch8_in;
  logic [86:0] zll_main_loop81_in;
  logic [86:0] zll_main_putins11_in;
  logic [69:0] zll_main_putins11_out;
  logic [69:0] zll_main_loop225_in;
  logic [142:0] zll_main_loop225_out;
  logic [142:0] zll_main_loop169_in;
  logic [142:0] zll_main_loop63_in;
  logic [69:0] zll_main_loop193_in;
  logic [69:0] main_incrpc_in;
  logic [69:0] main_incrpc_out;
  logic [69:0] zll_main_loop225_inR1;
  logic [142:0] zll_main_loop225_outR1;
  logic [142:0] zll_main_loop197_in;
  logic [142:0] zll_main_loop166_in;
  logic [69:0] zll_main_loop163_in;
  logic [69:0] main_getpc_in;
  logic [75:0] main_getpc_out;
  logic [75:0] zll_main_loop112_in;
  logic [69:0] zll_main_loop112_out;
  logic [69:0] zll_main_loop225_inR2;
  logic [142:0] zll_main_loop225_outR2;
  logic [142:0] zll_main_loop31_in;
  logic [142:0] zll_main_loop171_in;
  logic [69:0] zll_main_loop49_in;
  logic [69:0] main_getout_in;
  logic [84:0] main_getout_out;
  logic [84:0] zll_main_loop140_in;
  logic [142:0] zll_main_loop140_out;
  logic [142:0] zll_main_loop46_in;
  logic [142:0] zll_main_loop80_in;
  logic [84:0] zll_main_loop47_in;
  logic [90:0] zll_pure_dispatch3_in;
  logic [86:0] zll_main_loop86_in;
  logic [86:0] zll_main_putins11_inR1;
  logic [69:0] zll_main_putins11_outR1;
  logic [69:0] zll_main_loop225_inR3;
  logic [142:0] zll_main_loop225_outR3;
  logic [142:0] zll_main_loop5_in;
  logic [142:0] zll_main_loop19_in;
  logic [69:0] zll_main_loop113_in;
  logic [69:0] main_getdatain_in;
  logic [69:0] main_getins_in;
  logic [86:0] main_getins_out;
  logic [86:0] zll_main_getdatain1_in;
  logic [86:0] zll_main_getdatain2_in;
  logic [16:0] zll_main_datain_in;
  logic [16:0] zll_main_datain2_in;
  logic [77:0] zll_main_loop135_in;
  logic [77:0] main_putreg1_in;
  logic [89:0] zll_main_putreg27_in;
  logic [69:0] zll_main_putreg27_out;
  logic [69:0] zll_main_loop225_inR4;
  logic [142:0] zll_main_loop225_outR4;
  logic [142:0] zll_main_loop221_in;
  logic [142:0] zll_main_loop221_out;
  logic [90:0] zll_pure_dispatch_in;
  logic [86:0] zll_main_reset11_in;
  logic [86:0] zll_main_putins11_inR2;
  logic [69:0] zll_main_putins11_outR2;
  logic [69:0] zll_main_loop225_inR5;
  logic [142:0] zll_main_loop225_outR5;
  logic [142:0] zll_main_reset4_in;
  logic [142:0] zll_main_reset39_in;
  logic [69:0] zll_main_reset10_in;
  logic [69:0] main_getpc_inR1;
  logic [75:0] main_getpc_outR1;
  logic [75:0] zll_main_loop112_inR1;
  logic [69:0] zll_main_loop112_outR1;
  logic [69:0] zll_main_loop225_inR6;
  logic [142:0] zll_main_loop225_outR6;
  logic [142:0] zll_main_reset29_in;
  logic [142:0] zll_main_reset45_in;
  logic [69:0] zll_main_reset37_in;
  logic [69:0] main_getout_inR1;
  logic [84:0] main_getout_outR1;
  logic [84:0] zll_main_loop140_inR1;
  logic [142:0] zll_main_loop140_outR1;
  logic [142:0] zll_main_reset46_in;
  logic [142:0] zll_main_reset33_in;
  logic [84:0] zll_main_reset36_in;
  logic [90:0] zll_pure_dispatch7_inR2;
  logic [142:0] zll_pure_dispatch7_outR2;
  logic [90:0] zll_pure_dispatch7_inR3;
  logic [142:0] zll_pure_dispatch7_outR3;
  logic [90:0] zll_pure_dispatch2_in;
  logic [86:0] zll_main_loop213_in;
  logic [86:0] zll_main_putins11_inR3;
  logic [69:0] zll_main_putins11_outR3;
  logic [69:0] zll_main_loop225_inR7;
  logic [142:0] zll_main_loop225_outR7;
  logic [142:0] zll_main_loop181_in;
  logic [142:0] zll_main_loop129_in;
  logic [69:0] zll_main_loop20_in;
  logic [69:0] main_incrpc_inR1;
  logic [69:0] main_incrpc_outR1;
  logic [69:0] zll_main_loop225_inR8;
  logic [142:0] zll_main_loop225_outR8;
  logic [142:0] zll_main_loop226_in;
  logic [142:0] zll_main_loop216_in;
  logic [69:0] zll_main_loop148_in;
  logic [69:0] main_getpc_inR2;
  logic [75:0] main_getpc_outR2;
  logic [75:0] zll_main_loop112_inR2;
  logic [69:0] zll_main_loop112_outR2;
  logic [69:0] zll_main_loop225_inR9;
  logic [142:0] zll_main_loop225_outR9;
  logic [142:0] zll_main_loop110_in;
  logic [142:0] zll_main_loop105_in;
  logic [69:0] zll_main_loop25_in;
  logic [69:0] main_getout_inR2;
  logic [84:0] main_getout_outR2;
  logic [84:0] zll_main_loop140_inR2;
  logic [142:0] zll_main_loop140_outR2;
  logic [142:0] zll_main_loop92_in;
  logic [142:0] zll_main_loop2_in;
  logic [84:0] zll_main_loop24_in;
  logic [90:0] zll_pure_dispatch7_inR4;
  logic [142:0] zll_pure_dispatch7_outR4;
  logic [53:0] __padding;
  logic [3:0] __resumption_tag;
  logic [69:0] __st0;
  logic [3:0] __resumption_tag_next;
  logic [69:0] __st0_next;
  assign zll_pure_dispatch7_in = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch7  inst (zll_pure_dispatch7_in[90:74], zll_pure_dispatch7_in[69:0], zll_pure_dispatch7_out);
  assign zll_pure_dispatch7_inR1 = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch7  instR1 (zll_pure_dispatch7_inR1[90:74], zll_pure_dispatch7_inR1[69:0], zll_pure_dispatch7_outR1);
  assign zll_pure_dispatch8_in = {__in0, {__resumption_tag, __st0}};
  assign zll_main_loop81_in = {zll_pure_dispatch8_in[90:74], zll_pure_dispatch8_in[69:0]};
  assign zll_main_putins11_in = {zll_main_loop81_in[86:70], zll_main_loop81_in[69:0]};
  ZLL_Main_putIns11  instR2 (zll_main_putins11_in[86:70], zll_main_putins11_in[69:0], zll_main_putins11_out);
  assign zll_main_loop225_in = zll_main_putins11_out;
  ZLL_Main_loop225  instR3 (zll_main_loop225_in[69:0], zll_main_loop225_out);
  assign zll_main_loop169_in = zll_main_loop225_out;
  assign zll_main_loop63_in = zll_main_loop169_in[142:0];
  assign zll_main_loop193_in = zll_main_loop63_in[69:0];
  assign main_incrpc_in = zll_main_loop193_in[69:0];
  Main_incrPC  instR4 (main_incrpc_in[69:0], main_incrpc_out);
  assign zll_main_loop225_inR1 = main_incrpc_out;
  ZLL_Main_loop225  instR5 (zll_main_loop225_inR1[69:0], zll_main_loop225_outR1);
  assign zll_main_loop197_in = zll_main_loop225_outR1;
  assign zll_main_loop166_in = zll_main_loop197_in[142:0];
  assign zll_main_loop163_in = zll_main_loop166_in[69:0];
  assign main_getpc_in = zll_main_loop163_in[69:0];
  Main_getPC  instR6 (main_getpc_in[69:0], main_getpc_out);
  assign zll_main_loop112_in = main_getpc_out;
  ZLL_Main_loop112  instR7 (zll_main_loop112_in[75:0], zll_main_loop112_out);
  assign zll_main_loop225_inR2 = zll_main_loop112_out;
  ZLL_Main_loop225  instR8 (zll_main_loop225_inR2[69:0], zll_main_loop225_outR2);
  assign zll_main_loop31_in = zll_main_loop225_outR2;
  assign zll_main_loop171_in = zll_main_loop31_in[142:0];
  assign zll_main_loop49_in = zll_main_loop171_in[69:0];
  assign main_getout_in = zll_main_loop49_in[69:0];
  Main_getOut  instR9 (main_getout_in[69:0], main_getout_out);
  assign zll_main_loop140_in = main_getout_out;
  ZLL_Main_loop140  instR10 (zll_main_loop140_in[84:0], zll_main_loop140_out);
  assign zll_main_loop46_in = zll_main_loop140_out;
  assign zll_main_loop80_in = zll_main_loop46_in[142:0];
  assign zll_main_loop47_in = {zll_main_loop80_in[84:70], zll_main_loop80_in[69:0]};
  assign zll_pure_dispatch3_in = {__in0, {__resumption_tag, __st0}};
  assign zll_main_loop86_in = {zll_pure_dispatch3_in[90:74], zll_pure_dispatch3_in[69:0]};
  assign zll_main_putins11_inR1 = {zll_main_loop86_in[86:70], zll_main_loop86_in[69:0]};
  ZLL_Main_putIns11  instR11 (zll_main_putins11_inR1[86:70], zll_main_putins11_inR1[69:0], zll_main_putins11_outR1);
  assign zll_main_loop225_inR3 = zll_main_putins11_outR1;
  ZLL_Main_loop225  instR12 (zll_main_loop225_inR3[69:0], zll_main_loop225_outR3);
  assign zll_main_loop5_in = zll_main_loop225_outR3;
  assign zll_main_loop19_in = zll_main_loop5_in[142:0];
  assign zll_main_loop113_in = zll_main_loop19_in[69:0];
  assign main_getdatain_in = zll_main_loop113_in[69:0];
  assign main_getins_in = main_getdatain_in[69:0];
  Main_getIns  instR13 (main_getins_in[69:0], main_getins_out);
  assign zll_main_getdatain1_in = main_getins_out;
  assign zll_main_getdatain2_in = zll_main_getdatain1_in[86:0];
  assign zll_main_datain_in = zll_main_getdatain2_in[86:70];
  assign zll_main_datain2_in = zll_main_datain_in[16:0];
  assign zll_main_loop135_in = {zll_main_datain2_in[7:0], zll_main_getdatain2_in[69:0]};
  assign main_putreg1_in = zll_main_loop135_in[77:0];
  assign zll_main_putreg27_in = {main_putreg1_in[77:70], 4'h0, main_putreg1_in[77:70], main_putreg1_in[69:0]};
  ZLL_Main_putReg27  instR14 (zll_main_putreg27_in[89:82], zll_main_putreg27_in[81:80], zll_main_putreg27_in[79:70], zll_main_putreg27_in[69:0], zll_main_putreg27_out);
  assign zll_main_loop225_inR4 = zll_main_putreg27_out;
  ZLL_Main_loop225  instR15 (zll_main_loop225_inR4[69:0], zll_main_loop225_outR4);
  assign zll_main_loop221_in = zll_main_loop225_outR4;
  ZLL_Main_loop221  instR16 (zll_main_loop221_in[142:0], zll_main_loop221_out);
  assign zll_pure_dispatch_in = {__in0, {__resumption_tag, __st0}};
  assign zll_main_reset11_in = {zll_pure_dispatch_in[90:74], zll_pure_dispatch_in[69:0]};
  assign zll_main_putins11_inR2 = {zll_main_reset11_in[86:70], zll_main_reset11_in[69:0]};
  ZLL_Main_putIns11  instR17 (zll_main_putins11_inR2[86:70], zll_main_putins11_inR2[69:0], zll_main_putins11_outR2);
  assign zll_main_loop225_inR5 = zll_main_putins11_outR2;
  ZLL_Main_loop225  instR18 (zll_main_loop225_inR5[69:0], zll_main_loop225_outR5);
  assign zll_main_reset4_in = zll_main_loop225_outR5;
  assign zll_main_reset39_in = zll_main_reset4_in[142:0];
  assign zll_main_reset10_in = zll_main_reset39_in[69:0];
  assign main_getpc_inR1 = zll_main_reset10_in[69:0];
  Main_getPC  instR19 (main_getpc_inR1[69:0], main_getpc_outR1);
  assign zll_main_loop112_inR1 = main_getpc_outR1;
  ZLL_Main_loop112  instR20 (zll_main_loop112_inR1[75:0], zll_main_loop112_outR1);
  assign zll_main_loop225_inR6 = zll_main_loop112_outR1;
  ZLL_Main_loop225  instR21 (zll_main_loop225_inR6[69:0], zll_main_loop225_outR6);
  assign zll_main_reset29_in = zll_main_loop225_outR6;
  assign zll_main_reset45_in = zll_main_reset29_in[142:0];
  assign zll_main_reset37_in = zll_main_reset45_in[69:0];
  assign main_getout_inR1 = zll_main_reset37_in[69:0];
  Main_getOut  instR22 (main_getout_inR1[69:0], main_getout_outR1);
  assign zll_main_loop140_inR1 = main_getout_outR1;
  ZLL_Main_loop140  instR23 (zll_main_loop140_inR1[84:0], zll_main_loop140_outR1);
  assign zll_main_reset46_in = zll_main_loop140_outR1;
  assign zll_main_reset33_in = zll_main_reset46_in[142:0];
  assign zll_main_reset36_in = {zll_main_reset33_in[84:70], zll_main_reset33_in[69:0]};
  assign zll_pure_dispatch7_inR2 = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch7  instR24 (zll_pure_dispatch7_inR2[90:74], zll_pure_dispatch7_inR2[69:0], zll_pure_dispatch7_outR2);
  assign zll_pure_dispatch7_inR3 = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch7  instR25 (zll_pure_dispatch7_inR3[90:74], zll_pure_dispatch7_inR3[69:0], zll_pure_dispatch7_outR3);
  assign zll_pure_dispatch2_in = {__in0, {__resumption_tag, __st0}};
  assign zll_main_loop213_in = {zll_pure_dispatch2_in[90:74], zll_pure_dispatch2_in[69:0]};
  assign zll_main_putins11_inR3 = {zll_main_loop213_in[86:70], zll_main_loop213_in[69:0]};
  ZLL_Main_putIns11  instR26 (zll_main_putins11_inR3[86:70], zll_main_putins11_inR3[69:0], zll_main_putins11_outR3);
  assign zll_main_loop225_inR7 = zll_main_putins11_outR3;
  ZLL_Main_loop225  instR27 (zll_main_loop225_inR7[69:0], zll_main_loop225_outR7);
  assign zll_main_loop181_in = zll_main_loop225_outR7;
  assign zll_main_loop129_in = zll_main_loop181_in[142:0];
  assign zll_main_loop20_in = zll_main_loop129_in[69:0];
  assign main_incrpc_inR1 = zll_main_loop20_in[69:0];
  Main_incrPC  instR28 (main_incrpc_inR1[69:0], main_incrpc_outR1);
  assign zll_main_loop225_inR8 = main_incrpc_outR1;
  ZLL_Main_loop225  instR29 (zll_main_loop225_inR8[69:0], zll_main_loop225_outR8);
  assign zll_main_loop226_in = zll_main_loop225_outR8;
  assign zll_main_loop216_in = zll_main_loop226_in[142:0];
  assign zll_main_loop148_in = zll_main_loop216_in[69:0];
  assign main_getpc_inR2 = zll_main_loop148_in[69:0];
  Main_getPC  instR30 (main_getpc_inR2[69:0], main_getpc_outR2);
  assign zll_main_loop112_inR2 = main_getpc_outR2;
  ZLL_Main_loop112  instR31 (zll_main_loop112_inR2[75:0], zll_main_loop112_outR2);
  assign zll_main_loop225_inR9 = zll_main_loop112_outR2;
  ZLL_Main_loop225  instR32 (zll_main_loop225_inR9[69:0], zll_main_loop225_outR9);
  assign zll_main_loop110_in = zll_main_loop225_outR9;
  assign zll_main_loop105_in = zll_main_loop110_in[142:0];
  assign zll_main_loop25_in = zll_main_loop105_in[69:0];
  assign main_getout_inR2 = zll_main_loop25_in[69:0];
  Main_getOut  instR33 (main_getout_inR2[69:0], main_getout_outR2);
  assign zll_main_loop140_inR2 = main_getout_outR2;
  ZLL_Main_loop140  instR34 (zll_main_loop140_inR2[84:0], zll_main_loop140_outR2);
  assign zll_main_loop92_in = zll_main_loop140_outR2;
  assign zll_main_loop2_in = zll_main_loop92_in[142:0];
  assign zll_main_loop24_in = {zll_main_loop2_in[84:70], zll_main_loop2_in[69:0]};
  assign zll_pure_dispatch7_inR4 = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch7  instR35 (zll_pure_dispatch7_inR4[90:74], zll_pure_dispatch7_inR4[69:0], zll_pure_dispatch7_outR4);
  assign {__padding, __out0, __resumption_tag_next, __st0_next} = (zll_pure_dispatch7_inR4[73:70] == 4'h1) ? zll_pure_dispatch7_outR4 : ((zll_pure_dispatch2_in[73:70] == 4'h2) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop24_in[84:70], 4'h8, zll_main_loop24_in[69:0]} : ((zll_pure_dispatch7_inR3[73:70] == 4'h3) ? zll_pure_dispatch7_outR3 : ((zll_pure_dispatch7_inR2[73:70] == 4'h4) ? zll_pure_dispatch7_outR2 : ((zll_pure_dispatch_in[73:70] == 4'h5) ? {{1'h1, {6'h35{1'h0}}}, zll_main_reset36_in[84:70], 4'h1, zll_main_reset36_in[69:0]} : ((zll_pure_dispatch3_in[73:70] == 4'h6) ? zll_main_loop221_out : ((zll_pure_dispatch8_in[73:70] == 4'h7) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop47_in[84:70], 4'h6, zll_main_loop47_in[69:0]} : ((zll_pure_dispatch7_inR1[73:70] == 4'h8) ? zll_pure_dispatch7_outR1 : zll_pure_dispatch7_out)))))));
  initial {__resumption_tag, __st0} = {4'h5, {7'h46{1'h0}}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      {__resumption_tag, __st0} <= {4'h5, {7'h46{1'h0}}};
    end else begin
      {__resumption_tag, __st0} <= {__resumption_tag_next, __st0_next};
    end
  end
endmodule

module ZLL_Main_loop225 (input logic [69:0] arg0,
  output logic [142:0] res);
  assign res = {{2'h1, {7'h47{1'h0}}}, arg0};
endmodule

module ZLL_Main_r27 (input logic [7:0] arg0,
  input logic [7:0] arg1,
  input logic [5:0] arg2,
  input logic [16:0] arg3,
  input logic [14:0] arg4,
  output logic [7:0] res);
  logic [45:0] zll_main_r35_in;
  logic [7:0] zll_main_r35_out;
  assign zll_main_r35_in = {arg0, arg2, arg3, arg4};
  ZLL_Main_r35  inst (zll_main_r35_in[45:38], zll_main_r35_in[37:32], zll_main_r35_in[31:15], zll_main_r35_in[14:0], zll_main_r35_out);
  assign res = zll_main_r35_out;
endmodule

module ZLL_Main_loop221 (input logic [142:0] arg0,
  output logic [142:0] res);
  logic [142:0] zll_main_loop214_in;
  logic [69:0] main_loop_in;
  logic [69:0] main_getinstr_in;
  logic [69:0] main_getins_in;
  logic [86:0] main_getins_out;
  logic [86:0] zll_main_getinstr_in;
  logic [86:0] zll_main_getinstr1_in;
  logic [16:0] zll_main_instrin_in;
  logic [16:0] zll_main_instrin1_in;
  logic [78:0] zll_main_loop158_in;
  logic [78:0] zll_main_loop167_in;
  logic [142:0] zll_main_loop18_in;
  logic [142:0] zll_main_loop_in;
  logic [78:0] zll_main_loop211_in;
  logic [139:0] zll_main_loop73_in;
  logic [139:0] zll_main_loop121_in;
  logic [151:0] zll_main_loop58_in;
  logic [151:0] zll_main_loop223_in;
  logic [148:0] zll_main_loop215_in;
  logic [78:0] zll_main_loop199_in;
  logic [75:0] zll_main_loop50_in;
  logic [75:0] zll_main_loop52_in;
  logic [69:0] main_getreg1_in;
  logic [77:0] main_getreg1_out;
  logic [83:0] zll_main_loop222_in;
  logic [83:0] zll_main_bnz2_in;
  logic [15:0] binop_in;
  logic [84:0] zll_main_bnz4_in;
  logic [15:0] binop_inR1;
  logic [76:0] zll_main_bnz3_in;
  logic [76:0] zll_main_bnz6_in;
  logic [75:0] zll_main_bnz1_in;
  logic [75:0] zll_main_putpc14_in;
  logic [69:0] zll_main_putpc14_out;
  logic [70:0] zll_main_nand9_in;
  logic [69:0] main_incrpc_in;
  logic [69:0] main_incrpc_out;
  logic [69:0] zll_main_loop225_in;
  logic [142:0] zll_main_loop225_out;
  logic [142:0] zll_main_loop179_in;
  logic [142:0] zll_main_loop116_in;
  logic [69:0] zll_main_loop35_in;
  logic [69:0] main_getpc_in;
  logic [75:0] main_getpc_out;
  logic [75:0] zll_main_loop112_in;
  logic [69:0] zll_main_loop112_out;
  logic [69:0] zll_main_loop225_inR1;
  logic [142:0] zll_main_loop225_outR1;
  logic [142:0] zll_main_loop126_in;
  logic [142:0] zll_main_loop155_in;
  logic [69:0] zll_main_loop79_in;
  logic [69:0] main_getout_in;
  logic [84:0] main_getout_out;
  logic [84:0] zll_main_loop140_in;
  logic [142:0] zll_main_loop140_out;
  logic [142:0] zll_main_loop91_in;
  logic [142:0] zll_main_loop160_in;
  logic [84:0] zll_main_loop89_in;
  logic [78:0] zll_main_loop187_in;
  logic [75:0] zll_main_loop32_in;
  logic [75:0] zll_main_loop101_in;
  logic [75:0] zll_main_loop99_in;
  logic [71:0] main_getreg_in;
  logic [77:0] main_getreg_out;
  logic [81:0] zll_main_loop127_in;
  logic [81:0] zll_main_loop68_in;
  logic [81:0] zll_main_loop87_in;
  logic [81:0] zll_main_nand4_in;
  logic [71:0] main_getreg_inR1;
  logic [77:0] main_getreg_outR1;
  logic [87:0] zll_main_nand5_in;
  logic [87:0] zll_main_nand3_in;
  logic [15:0] binop_inR2;
  logic [7:0] unop_in;
  logic [79:0] main_putreg_in;
  logic [89:0] zll_main_putreg27_in;
  logic [69:0] zll_main_putreg27_out;
  logic [69:0] main_incrpc_inR1;
  logic [69:0] main_incrpc_outR1;
  logic [69:0] zll_main_loop225_inR2;
  logic [142:0] zll_main_loop225_outR2;
  logic [142:0] zll_main_loop88_in;
  logic [142:0] zll_main_loop84_in;
  logic [69:0] zll_main_loop15_in;
  logic [69:0] main_getpc_inR1;
  logic [75:0] main_getpc_outR1;
  logic [75:0] zll_main_loop112_inR1;
  logic [69:0] zll_main_loop112_outR1;
  logic [69:0] zll_main_loop225_inR3;
  logic [142:0] zll_main_loop225_outR3;
  logic [142:0] zll_main_loop118_in;
  logic [142:0] zll_main_loop204_in;
  logic [69:0] zll_main_loop178_in;
  logic [69:0] main_getout_inR1;
  logic [84:0] main_getout_outR1;
  logic [84:0] zll_main_loop140_inR1;
  logic [142:0] zll_main_loop140_outR1;
  logic [142:0] zll_main_loop30_in;
  logic [142:0] zll_main_loop201_in;
  logic [84:0] zll_main_loop209_in;
  logic [78:0] zll_main_loop71_in;
  logic [75:0] zll_main_loop95_in;
  logic [75:0] zll_main_loop82_in;
  logic [69:0] main_getreg1_inR1;
  logic [77:0] main_getreg1_outR1;
  logic [83:0] zll_main_loop132_in;
  logic [83:0] zll_main_st_in;
  logic [75:0] zll_main_putaddrout1_in;
  logic [69:0] zll_main_putaddrout1_out;
  logic [77:0] zll_main_st3_in;
  logic [77:0] zll_main_putdataout3_in;
  logic [69:0] main_getout_inR2;
  logic [84:0] main_getout_outR2;
  logic [92:0] zll_main_putdataout4_in;
  logic [92:0] zll_main_putdataout7_in;
  logic [22:0] zll_main_putdataout6_in;
  logic [22:0] zll_main_putdataout11_in;
  logic [22:0] zll_main_putdataout_in;
  logic [84:0] zll_main_putout5_in;
  logic [69:0] zll_main_putout5_out;
  logic [69:0] main_putweout1_in;
  logic [70:0] zll_main_putweout2_in;
  logic [69:0] zll_main_putweout2_out;
  logic [69:0] zll_main_loop225_inR4;
  logic [142:0] zll_main_loop225_outR4;
  logic [142:0] zll_main_loop159_in;
  logic [142:0] zll_main_loop38_in;
  logic [69:0] zll_main_loop14_in;
  logic [69:0] main_getout_inR3;
  logic [84:0] main_getout_outR3;
  logic [84:0] zll_main_loop140_inR2;
  logic [142:0] zll_main_loop140_outR2;
  logic [142:0] zll_main_loop104_in;
  logic [142:0] zll_main_loop78_in;
  logic [84:0] zll_main_loop41_in;
  logic [78:0] zll_main_loop100_in;
  logic [75:0] zll_main_loop180_in;
  logic [75:0] zll_main_loop142_in;
  logic [75:0] zll_main_putaddrout1_inR1;
  logic [69:0] zll_main_putaddrout1_outR1;
  logic [69:0] main_putweout_in;
  logic [69:0] main_putweout_out;
  logic [69:0] zll_main_loop225_inR5;
  logic [142:0] zll_main_loop225_outR5;
  logic [142:0] zll_main_loop173_in;
  logic [142:0] zll_main_loop65_in;
  logic [69:0] zll_main_loop123_in;
  logic [69:0] main_getout_inR4;
  logic [84:0] main_getout_outR4;
  logic [84:0] zll_main_loop140_inR3;
  logic [142:0] zll_main_loop140_outR3;
  logic [142:0] zll_main_loop128_in;
  logic [142:0] zll_main_loop10_in;
  logic [84:0] zll_main_loop21_in;
  logic [78:0] zll_main_loop9_in;
  logic [69:0] zll_main_loop76_in;
  logic [69:0] main_incrpc_inR2;
  logic [69:0] main_incrpc_outR2;
  logic [69:0] zll_main_loop225_inR6;
  logic [142:0] zll_main_loop225_outR6;
  logic [142:0] zll_main_loop147_in;
  logic [142:0] zll_main_loop106_in;
  logic [69:0] zll_main_loop124_in;
  logic [69:0] main_getpc_inR2;
  logic [75:0] main_getpc_outR2;
  logic [75:0] zll_main_loop112_inR2;
  logic [69:0] zll_main_loop112_outR2;
  logic [69:0] zll_main_loop225_inR7;
  logic [142:0] zll_main_loop225_outR7;
  logic [142:0] zll_main_loop217_in;
  logic [142:0] zll_main_loop138_in;
  logic [69:0] zll_main_loop139_in;
  logic [69:0] main_getout_inR5;
  logic [84:0] main_getout_outR5;
  logic [84:0] zll_main_loop140_inR4;
  logic [142:0] zll_main_loop140_outR4;
  logic [142:0] zll_main_loop13_in;
  logic [142:0] zll_main_loop198_in;
  logic [84:0] zll_main_loop200_in;
  assign zll_main_loop214_in = arg0;
  assign main_loop_in = zll_main_loop214_in[69:0];
  assign main_getinstr_in = main_loop_in[69:0];
  assign main_getins_in = main_getinstr_in[69:0];
  Main_getIns  inst (main_getins_in[69:0], main_getins_out);
  assign zll_main_getinstr_in = main_getins_out;
  assign zll_main_getinstr1_in = zll_main_getinstr_in[86:0];
  assign zll_main_instrin_in = zll_main_getinstr1_in[86:70];
  assign zll_main_instrin1_in = zll_main_instrin_in[16:0];
  assign zll_main_loop158_in = {zll_main_instrin1_in[16:8], zll_main_getinstr1_in[69:0]};
  assign zll_main_loop167_in = zll_main_loop158_in[78:0];
  assign zll_main_loop18_in = {{7'h40{1'h0}}, zll_main_loop167_in[78:70], zll_main_loop167_in[69:0]};
  assign zll_main_loop_in = zll_main_loop18_in[142:0];
  assign zll_main_loop211_in = {zll_main_loop_in[78:70], zll_main_loop_in[69:0]};
  assign zll_main_loop73_in = {zll_main_loop211_in[69:0], zll_main_loop211_in[69:0]};
  assign zll_main_loop121_in = zll_main_loop73_in[139:0];
  assign zll_main_loop58_in = {zll_main_loop211_in[78:70], {3'h3, zll_main_loop121_in[139:70], zll_main_loop121_in[69:0]}};
  assign zll_main_loop223_in = {zll_main_loop58_in[151:143], zll_main_loop58_in[142:0]};
  assign zll_main_loop215_in = {zll_main_loop223_in[151:143], zll_main_loop223_in[139:70], zll_main_loop223_in[69:0]};
  assign zll_main_loop199_in = {zll_main_loop215_in[69:0], zll_main_loop215_in[148:140]};
  assign zll_main_loop50_in = {zll_main_loop199_in[78:9], zll_main_loop199_in[5:0]};
  assign zll_main_loop52_in = {zll_main_loop50_in[5:0], zll_main_loop50_in[75:6]};
  assign main_getreg1_in = zll_main_loop52_in[69:0];
  Main_getReg1  instR1 (main_getreg1_in[69:0], main_getreg1_out);
  assign zll_main_loop222_in = {zll_main_loop52_in[75:70], main_getreg1_out};
  assign zll_main_bnz2_in = {zll_main_loop222_in[83:78], zll_main_loop222_in[77:0]};
  assign binop_in = {zll_main_bnz2_in[77:70], 8'h0};
  assign zll_main_bnz4_in = {zll_main_bnz2_in[77:70], zll_main_bnz2_in[83:78], binop_in[15:8] == binop_in[7:0], zll_main_bnz2_in[69:0]};
  assign binop_inR1 = {zll_main_bnz4_in[84:77], 8'h0};
  assign zll_main_bnz3_in = {zll_main_bnz4_in[76:71], binop_inR1[15:8] == binop_inR1[7:0], zll_main_bnz4_in[69:0]};
  assign zll_main_bnz6_in = {zll_main_bnz3_in[69:0], zll_main_bnz3_in[76:71], zll_main_bnz3_in[70]};
  assign zll_main_bnz1_in = {zll_main_bnz6_in[76:7], zll_main_bnz6_in[6:1]};
  assign zll_main_putpc14_in = {zll_main_bnz1_in[5:0], zll_main_bnz1_in[75:6]};
  ZLL_Main_putPC14  instR2 (zll_main_putpc14_in[75:70], zll_main_putpc14_in[69:0], zll_main_putpc14_out);
  assign zll_main_nand9_in = {zll_main_bnz4_in[69:0], zll_main_bnz4_in[70]};
  assign main_incrpc_in = zll_main_nand9_in[70:1];
  Main_incrPC  instR3 (main_incrpc_in[69:0], main_incrpc_out);
  assign zll_main_loop225_in = (zll_main_nand9_in[0] == 1'h1) ? main_incrpc_out : zll_main_putpc14_out;
  ZLL_Main_loop225  instR4 (zll_main_loop225_in[69:0], zll_main_loop225_out);
  assign zll_main_loop179_in = zll_main_loop225_out;
  assign zll_main_loop116_in = zll_main_loop179_in[142:0];
  assign zll_main_loop35_in = zll_main_loop116_in[69:0];
  assign main_getpc_in = zll_main_loop35_in[69:0];
  Main_getPC  instR5 (main_getpc_in[69:0], main_getpc_out);
  assign zll_main_loop112_in = main_getpc_out;
  ZLL_Main_loop112  instR6 (zll_main_loop112_in[75:0], zll_main_loop112_out);
  assign zll_main_loop225_inR1 = zll_main_loop112_out;
  ZLL_Main_loop225  instR7 (zll_main_loop225_inR1[69:0], zll_main_loop225_outR1);
  assign zll_main_loop126_in = zll_main_loop225_outR1;
  assign zll_main_loop155_in = zll_main_loop126_in[142:0];
  assign zll_main_loop79_in = zll_main_loop155_in[69:0];
  assign main_getout_in = zll_main_loop79_in[69:0];
  Main_getOut  instR8 (main_getout_in[69:0], main_getout_out);
  assign zll_main_loop140_in = main_getout_out;
  ZLL_Main_loop140  instR9 (zll_main_loop140_in[84:0], zll_main_loop140_out);
  assign zll_main_loop91_in = zll_main_loop140_out;
  assign zll_main_loop160_in = zll_main_loop91_in[142:0];
  assign zll_main_loop89_in = {zll_main_loop160_in[84:70], zll_main_loop160_in[69:0]};
  assign zll_main_loop187_in = {zll_main_loop215_in[69:0], zll_main_loop215_in[148:140]};
  assign zll_main_loop32_in = {zll_main_loop187_in[78:9], zll_main_loop187_in[5:4], zll_main_loop187_in[3:2], zll_main_loop187_in[1:0]};
  assign zll_main_loop101_in = {zll_main_loop32_in[5:4], zll_main_loop32_in[75:6], zll_main_loop32_in[3:2], zll_main_loop32_in[1:0]};
  assign zll_main_loop99_in = {zll_main_loop101_in[75:74], zll_main_loop101_in[3:2], zll_main_loop101_in[1:0], zll_main_loop101_in[73:4]};
  assign main_getreg_in = {zll_main_loop99_in[73:72], zll_main_loop99_in[69:0]};
  Main_getReg  instR10 (main_getreg_in[71:70], main_getreg_in[69:0], main_getreg_out);
  assign zll_main_loop127_in = {zll_main_loop99_in[71:70], zll_main_loop99_in[75:74], main_getreg_out};
  assign zll_main_loop68_in = {zll_main_loop127_in[81:80], zll_main_loop127_in[79:78], zll_main_loop127_in[77:0]};
  assign zll_main_loop87_in = {zll_main_loop68_in[79:78], zll_main_loop68_in[81:80], zll_main_loop68_in[77:70], zll_main_loop68_in[69:0]};
  assign zll_main_nand4_in = {zll_main_loop87_in[79:78], zll_main_loop87_in[81:80], zll_main_loop87_in[77:70], zll_main_loop87_in[69:0]};
  assign main_getreg_inR1 = {zll_main_nand4_in[81:80], zll_main_nand4_in[69:0]};
  Main_getReg  instR11 (main_getreg_inR1[71:70], main_getreg_inR1[69:0], main_getreg_outR1);
  assign zll_main_nand5_in = {zll_main_nand4_in[77:70], zll_main_nand4_in[79:78], main_getreg_outR1};
  assign zll_main_nand3_in = {zll_main_nand5_in[87:80], zll_main_nand5_in[79:78], zll_main_nand5_in[77:0]};
  assign binop_inR2 = {zll_main_nand3_in[87:80], zll_main_nand3_in[77:70]};
  assign unop_in = binop_inR2[15:8] & binop_inR2[7:0];
  assign main_putreg_in = {zll_main_nand3_in[79:78], ~unop_in[7:0], zll_main_nand3_in[69:0]};
  assign zll_main_putreg27_in = {main_putreg_in[77:70], main_putreg_in[79:78], main_putreg_in[79:78], main_putreg_in[77:70], main_putreg_in[69:0]};
  ZLL_Main_putReg27  instR12 (zll_main_putreg27_in[89:82], zll_main_putreg27_in[81:80], zll_main_putreg27_in[79:70], zll_main_putreg27_in[69:0], zll_main_putreg27_out);
  assign main_incrpc_inR1 = zll_main_putreg27_out;
  Main_incrPC  instR13 (main_incrpc_inR1[69:0], main_incrpc_outR1);
  assign zll_main_loop225_inR2 = main_incrpc_outR1;
  ZLL_Main_loop225  instR14 (zll_main_loop225_inR2[69:0], zll_main_loop225_outR2);
  assign zll_main_loop88_in = zll_main_loop225_outR2;
  assign zll_main_loop84_in = zll_main_loop88_in[142:0];
  assign zll_main_loop15_in = zll_main_loop84_in[69:0];
  assign main_getpc_inR1 = zll_main_loop15_in[69:0];
  Main_getPC  instR15 (main_getpc_inR1[69:0], main_getpc_outR1);
  assign zll_main_loop112_inR1 = main_getpc_outR1;
  ZLL_Main_loop112  instR16 (zll_main_loop112_inR1[75:0], zll_main_loop112_outR1);
  assign zll_main_loop225_inR3 = zll_main_loop112_outR1;
  ZLL_Main_loop225  instR17 (zll_main_loop225_inR3[69:0], zll_main_loop225_outR3);
  assign zll_main_loop118_in = zll_main_loop225_outR3;
  assign zll_main_loop204_in = zll_main_loop118_in[142:0];
  assign zll_main_loop178_in = zll_main_loop204_in[69:0];
  assign main_getout_inR1 = zll_main_loop178_in[69:0];
  Main_getOut  instR18 (main_getout_inR1[69:0], main_getout_outR1);
  assign zll_main_loop140_inR1 = main_getout_outR1;
  ZLL_Main_loop140  instR19 (zll_main_loop140_inR1[84:0], zll_main_loop140_outR1);
  assign zll_main_loop30_in = zll_main_loop140_outR1;
  assign zll_main_loop201_in = zll_main_loop30_in[142:0];
  assign zll_main_loop209_in = {zll_main_loop201_in[84:70], zll_main_loop201_in[69:0]};
  assign zll_main_loop71_in = {zll_main_loop215_in[69:0], zll_main_loop215_in[148:140]};
  assign zll_main_loop95_in = {zll_main_loop71_in[78:9], zll_main_loop71_in[5:0]};
  assign zll_main_loop82_in = {zll_main_loop95_in[5:0], zll_main_loop95_in[75:6]};
  assign main_getreg1_inR1 = zll_main_loop82_in[69:0];
  Main_getReg1  instR20 (main_getreg1_inR1[69:0], main_getreg1_outR1);
  assign zll_main_loop132_in = {zll_main_loop82_in[75:70], main_getreg1_outR1};
  assign zll_main_st_in = {zll_main_loop132_in[83:78], zll_main_loop132_in[77:0]};
  assign zll_main_putaddrout1_in = {zll_main_st_in[83:78], zll_main_st_in[69:0]};
  ZLL_Main_putAddrOut1  instR21 (zll_main_putaddrout1_in[75:70], zll_main_putaddrout1_in[69:0], zll_main_putaddrout1_out);
  assign zll_main_st3_in = {zll_main_st_in[77:70], zll_main_putaddrout1_out};
  assign zll_main_putdataout3_in = {zll_main_st3_in[77:70], zll_main_st3_in[69:0]};
  assign main_getout_inR2 = zll_main_putdataout3_in[69:0];
  Main_getOut  instR22 (main_getout_inR2[69:0], main_getout_outR2);
  assign zll_main_putdataout4_in = {zll_main_putdataout3_in[77:70], main_getout_outR2};
  assign zll_main_putdataout7_in = {zll_main_putdataout4_in[92:85], zll_main_putdataout4_in[84:0]};
  assign zll_main_putdataout6_in = {zll_main_putdataout7_in[92:85], zll_main_putdataout7_in[84:70]};
  assign zll_main_putdataout11_in = {zll_main_putdataout6_in[22:15], zll_main_putdataout6_in[14:0]};
  assign zll_main_putdataout_in = {zll_main_putdataout11_in[22:15], zll_main_putdataout11_in[13:8], zll_main_putdataout11_in[14], zll_main_putdataout11_in[7:0]};
  assign zll_main_putout5_in = {{zll_main_putdataout_in[8], zll_main_putdataout_in[14:9], zll_main_putdataout_in[22:15]}, zll_main_putdataout7_in[69:0]};
  ZLL_Main_putOut5  instR23 (zll_main_putout5_in[84:70], zll_main_putout5_in[69:0], zll_main_putout5_out);
  assign main_putweout1_in = zll_main_putout5_out;
  assign zll_main_putweout2_in = {1'h1, main_putweout1_in[69:0]};
  ZLL_Main_putWeOut2  instR24 (zll_main_putweout2_in[70], zll_main_putweout2_in[69:0], zll_main_putweout2_out);
  assign zll_main_loop225_inR4 = zll_main_putweout2_out;
  ZLL_Main_loop225  instR25 (zll_main_loop225_inR4[69:0], zll_main_loop225_outR4);
  assign zll_main_loop159_in = zll_main_loop225_outR4;
  assign zll_main_loop38_in = zll_main_loop159_in[142:0];
  assign zll_main_loop14_in = zll_main_loop38_in[69:0];
  assign main_getout_inR3 = zll_main_loop14_in[69:0];
  Main_getOut  instR26 (main_getout_inR3[69:0], main_getout_outR3);
  assign zll_main_loop140_inR2 = main_getout_outR3;
  ZLL_Main_loop140  instR27 (zll_main_loop140_inR2[84:0], zll_main_loop140_outR2);
  assign zll_main_loop104_in = zll_main_loop140_outR2;
  assign zll_main_loop78_in = zll_main_loop104_in[142:0];
  assign zll_main_loop41_in = {zll_main_loop78_in[84:70], zll_main_loop78_in[69:0]};
  assign zll_main_loop100_in = {zll_main_loop215_in[69:0], zll_main_loop215_in[148:140]};
  assign zll_main_loop180_in = {zll_main_loop100_in[78:9], zll_main_loop100_in[5:0]};
  assign zll_main_loop142_in = {zll_main_loop180_in[5:0], zll_main_loop180_in[75:6]};
  assign zll_main_putaddrout1_inR1 = {zll_main_loop142_in[75:70], zll_main_loop142_in[69:0]};
  ZLL_Main_putAddrOut1  instR28 (zll_main_putaddrout1_inR1[75:70], zll_main_putaddrout1_inR1[69:0], zll_main_putaddrout1_outR1);
  assign main_putweout_in = zll_main_putaddrout1_outR1;
  Main_putWeOut  instR29 (main_putweout_in[69:0], main_putweout_out);
  assign zll_main_loop225_inR5 = main_putweout_out;
  ZLL_Main_loop225  instR30 (zll_main_loop225_inR5[69:0], zll_main_loop225_outR5);
  assign zll_main_loop173_in = zll_main_loop225_outR5;
  assign zll_main_loop65_in = zll_main_loop173_in[142:0];
  assign zll_main_loop123_in = zll_main_loop65_in[69:0];
  assign main_getout_inR4 = zll_main_loop123_in[69:0];
  Main_getOut  instR31 (main_getout_inR4[69:0], main_getout_outR4);
  assign zll_main_loop140_inR3 = main_getout_outR4;
  ZLL_Main_loop140  instR32 (zll_main_loop140_inR3[84:0], zll_main_loop140_outR3);
  assign zll_main_loop128_in = zll_main_loop140_outR3;
  assign zll_main_loop10_in = zll_main_loop128_in[142:0];
  assign zll_main_loop21_in = {zll_main_loop10_in[84:70], zll_main_loop10_in[69:0]};
  assign zll_main_loop9_in = {zll_main_loop215_in[69:0], zll_main_loop215_in[148:140]};
  assign zll_main_loop76_in = zll_main_loop9_in[78:9];
  assign main_incrpc_inR2 = zll_main_loop76_in[69:0];
  Main_incrPC  instR33 (main_incrpc_inR2[69:0], main_incrpc_outR2);
  assign zll_main_loop225_inR6 = main_incrpc_outR2;
  ZLL_Main_loop225  instR34 (zll_main_loop225_inR6[69:0], zll_main_loop225_outR6);
  assign zll_main_loop147_in = zll_main_loop225_outR6;
  assign zll_main_loop106_in = zll_main_loop147_in[142:0];
  assign zll_main_loop124_in = zll_main_loop106_in[69:0];
  assign main_getpc_inR2 = zll_main_loop124_in[69:0];
  Main_getPC  instR35 (main_getpc_inR2[69:0], main_getpc_outR2);
  assign zll_main_loop112_inR2 = main_getpc_outR2;
  ZLL_Main_loop112  instR36 (zll_main_loop112_inR2[75:0], zll_main_loop112_outR2);
  assign zll_main_loop225_inR7 = zll_main_loop112_outR2;
  ZLL_Main_loop225  instR37 (zll_main_loop225_inR7[69:0], zll_main_loop225_outR7);
  assign zll_main_loop217_in = zll_main_loop225_outR7;
  assign zll_main_loop138_in = zll_main_loop217_in[142:0];
  assign zll_main_loop139_in = zll_main_loop138_in[69:0];
  assign main_getout_inR5 = zll_main_loop139_in[69:0];
  Main_getOut  instR38 (main_getout_inR5[69:0], main_getout_outR5);
  assign zll_main_loop140_inR4 = main_getout_outR5;
  ZLL_Main_loop140  instR39 (zll_main_loop140_inR4[84:0], zll_main_loop140_outR4);
  assign zll_main_loop13_in = zll_main_loop140_outR4;
  assign zll_main_loop198_in = zll_main_loop13_in[142:0];
  assign zll_main_loop200_in = {zll_main_loop198_in[84:70], zll_main_loop198_in[69:0]};
  assign res = (zll_main_loop9_in[8:6] == 3'h0) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop200_in[84:70], 4'h0, zll_main_loop200_in[69:0]} : ((zll_main_loop100_in[8:6] == 3'h1) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop21_in[84:70], 4'h7, zll_main_loop21_in[69:0]} : ((zll_main_loop71_in[8:6] == 3'h2) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop41_in[84:70], 4'h2, zll_main_loop41_in[69:0]} : ((zll_main_loop187_in[8:6] == 3'h3) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop209_in[84:70], 4'h4, zll_main_loop209_in[69:0]} : {{1'h1, {6'h35{1'h0}}}, zll_main_loop89_in[84:70], 4'h3, zll_main_loop89_in[69:0]})));
endmodule

module ZLL_Main_putPC14 (input logic [5:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [145:0] zll_main_putpc11_in;
  logic [145:0] zll_main_putpc10_in;
  logic [75:0] zll_main_putpc13_in;
  logic [75:0] zll_main_putpc8_in;
  logic [75:0] zll_main_putpc6_in;
  logic [75:0] zll_main_putpc12_in;
  logic [69:0] zll_main_putpc7_in;
  assign zll_main_putpc11_in = {arg0, arg1, arg1};
  assign zll_main_putpc10_in = {zll_main_putpc11_in[145:140], zll_main_putpc11_in[139:0]};
  assign zll_main_putpc13_in = {zll_main_putpc10_in[145:140], zll_main_putpc10_in[139:70]};
  assign zll_main_putpc8_in = {zll_main_putpc13_in[75:70], zll_main_putpc13_in[69:0]};
  assign zll_main_putpc6_in = {zll_main_putpc8_in[75:70], zll_main_putpc8_in[53:46], zll_main_putpc8_in[69:62], zll_main_putpc8_in[61:54], zll_main_putpc8_in[45:38], zll_main_putpc8_in[37:32], zll_main_putpc8_in[31:15], zll_main_putpc8_in[14:0]};
  assign zll_main_putpc12_in = {zll_main_putpc6_in[75:70], zll_main_putpc6_in[45:38], zll_main_putpc6_in[69:62], zll_main_putpc6_in[61:54], zll_main_putpc6_in[53:46], zll_main_putpc6_in[37:32], zll_main_putpc6_in[31:15], zll_main_putpc6_in[14:0]};
  assign zll_main_putpc7_in = {zll_main_putpc12_in[75:70], zll_main_putpc12_in[69:62], zll_main_putpc12_in[61:54], zll_main_putpc12_in[53:46], zll_main_putpc12_in[45:38], zll_main_putpc12_in[31:15], zll_main_putpc12_in[14:0]};
  assign res = {zll_main_putpc7_in[47:40], zll_main_putpc7_in[39:32], zll_main_putpc7_in[55:48], zll_main_putpc7_in[63:56], zll_main_putpc7_in[69:64], zll_main_putpc7_in[31:15], zll_main_putpc7_in[14:0]};
endmodule

module Main_getReg1 (input logic [69:0] arg0,
  output logic [77:0] res);
  logic [73:0] zll_main_getreg6_in;
  logic [77:0] zll_main_getreg6_out;
  assign zll_main_getreg6_in = {4'h0, arg0};
  ZLL_Main_getReg6  inst (zll_main_getreg6_in[73:72], zll_main_getreg6_in[71:70], zll_main_getreg6_in[69:0], zll_main_getreg6_out);
  assign res = zll_main_getreg6_out;
endmodule

module ZLL_Pure_dispatch7 (input logic [16:0] arg0,
  input logic [69:0] arg1,
  output logic [142:0] res);
  logic [86:0] zll_main_loop220_in;
  logic [86:0] zll_main_putins11_in;
  logic [69:0] zll_main_putins11_out;
  logic [69:0] zll_main_loop225_in;
  logic [142:0] zll_main_loop225_out;
  logic [142:0] zll_main_loop221_in;
  logic [142:0] zll_main_loop221_out;
  assign zll_main_loop220_in = {arg0, arg1};
  assign zll_main_putins11_in = {zll_main_loop220_in[86:70], zll_main_loop220_in[69:0]};
  ZLL_Main_putIns11  inst (zll_main_putins11_in[86:70], zll_main_putins11_in[69:0], zll_main_putins11_out);
  assign zll_main_loop225_in = zll_main_putins11_out;
  ZLL_Main_loop225  instR1 (zll_main_loop225_in[69:0], zll_main_loop225_out);
  assign zll_main_loop221_in = zll_main_loop225_out;
  ZLL_Main_loop221  instR2 (zll_main_loop221_in[142:0], zll_main_loop221_out);
  assign res = zll_main_loop221_out;
endmodule

module Main_getReg (input logic [1:0] arg0,
  input logic [69:0] arg1,
  output logic [77:0] res);
  logic [73:0] zll_main_getreg6_in;
  logic [77:0] zll_main_getreg6_out;
  assign zll_main_getreg6_in = {arg0, arg0, arg1};
  ZLL_Main_getReg6  inst (zll_main_getreg6_in[73:72], zll_main_getreg6_in[71:70], zll_main_getreg6_in[69:0], zll_main_getreg6_out);
  assign res = zll_main_getreg6_out;
endmodule

module ZLL_Main_r35 (input logic [7:0] arg0,
  input logic [5:0] arg1,
  input logic [16:0] arg2,
  input logic [14:0] arg3,
  output logic [7:0] res);
  logic [39:0] zll_main_r25_in;
  logic [22:0] zll_main_r26_in;
  assign zll_main_r25_in = {arg0, arg2, arg3};
  assign zll_main_r26_in = {zll_main_r25_in[39:32], zll_main_r25_in[14:0]};
  assign res = zll_main_r26_in[22:15];
endmodule

module ZLL_Main_putIns11 (input logic [16:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [156:0] zll_main_putins12_in;
  logic [156:0] zll_main_putins1_in;
  logic [86:0] zll_main_putins2_in;
  logic [86:0] zll_main_putins3_in;
  logic [86:0] zll_main_putins4_in;
  logic [86:0] zll_main_putins9_in;
  logic [86:0] zll_main_putins14_in;
  assign zll_main_putins12_in = {arg0, arg1, arg1};
  assign zll_main_putins1_in = {zll_main_putins12_in[156:140], zll_main_putins12_in[139:0]};
  assign zll_main_putins2_in = {zll_main_putins1_in[156:140], zll_main_putins1_in[139:70]};
  assign zll_main_putins3_in = {zll_main_putins2_in[86:70], zll_main_putins2_in[69:0]};
  assign zll_main_putins4_in = {zll_main_putins3_in[86:70], zll_main_putins3_in[53:46], zll_main_putins3_in[69:62], zll_main_putins3_in[61:54], zll_main_putins3_in[45:38], zll_main_putins3_in[37:32], zll_main_putins3_in[31:15], zll_main_putins3_in[14:0]};
  assign zll_main_putins9_in = {zll_main_putins4_in[86:70], zll_main_putins4_in[45:38], zll_main_putins4_in[69:62], zll_main_putins4_in[61:54], zll_main_putins4_in[53:46], zll_main_putins4_in[37:32], zll_main_putins4_in[31:15], zll_main_putins4_in[14:0]};
  assign zll_main_putins14_in = {zll_main_putins9_in[86:70], zll_main_putins9_in[69:62], zll_main_putins9_in[37:32], zll_main_putins9_in[61:54], zll_main_putins9_in[53:46], zll_main_putins9_in[45:38], zll_main_putins9_in[31:15], zll_main_putins9_in[14:0]};
  assign res = {zll_main_putins14_in[47:40], zll_main_putins14_in[39:32], zll_main_putins14_in[55:48], zll_main_putins14_in[69:62], zll_main_putins14_in[61:56], zll_main_putins14_in[86:70], zll_main_putins14_in[14:0]};
endmodule

module ZLL_Main_loop140 (input logic [84:0] arg0,
  output logic [142:0] res);
  logic [84:0] zll_main_loop207_in;
  assign zll_main_loop207_in = arg0;
  assign res = {{3'h1, {6'h37{1'h0}}}, zll_main_loop207_in[84:70], zll_main_loop207_in[69:0]};
endmodule

module Main_getIns (input logic [69:0] arg0,
  output logic [86:0] res);
  logic [139:0] zll_main_getins2_in;
  logic [139:0] zll_main_getins1_in;
  logic [69:0] zll_main_inputs5_in;
  logic [69:0] zll_main_inputs7_in;
  logic [61:0] zll_main_inputs6_in;
  logic [53:0] zll_main_inputs4_in;
  logic [45:0] zll_main_inputs_in;
  logic [37:0] zll_main_inputs1_in;
  logic [31:0] zll_main_inputs2_in;
  assign zll_main_getins2_in = {arg0, arg0};
  assign zll_main_getins1_in = zll_main_getins2_in[139:0];
  assign zll_main_inputs5_in = zll_main_getins1_in[139:70];
  assign zll_main_inputs7_in = zll_main_inputs5_in[69:0];
  assign zll_main_inputs6_in = {zll_main_inputs7_in[61:54], zll_main_inputs7_in[53:46], zll_main_inputs7_in[45:38], zll_main_inputs7_in[37:32], zll_main_inputs7_in[31:15], zll_main_inputs7_in[14:0]};
  assign zll_main_inputs4_in = {zll_main_inputs6_in[53:46], zll_main_inputs6_in[45:38], zll_main_inputs6_in[37:32], zll_main_inputs6_in[31:15], zll_main_inputs6_in[14:0]};
  assign zll_main_inputs_in = {zll_main_inputs4_in[45:38], zll_main_inputs4_in[37:32], zll_main_inputs4_in[31:15], zll_main_inputs4_in[14:0]};
  assign zll_main_inputs1_in = {zll_main_inputs_in[37:32], zll_main_inputs_in[31:15], zll_main_inputs_in[14:0]};
  assign zll_main_inputs2_in = {zll_main_inputs1_in[31:15], zll_main_inputs1_in[14:0]};
  assign res = {zll_main_inputs2_in[31:15], zll_main_getins1_in[69:0]};
endmodule

module ZLL_Main_loop112 (input logic [75:0] arg0,
  output logic [69:0] res);
  logic [75:0] zll_main_finishinstr1_in;
  logic [75:0] zll_main_putaddrout1_in;
  logic [69:0] zll_main_putaddrout1_out;
  logic [69:0] main_putweout_in;
  logic [69:0] main_putweout_out;
  assign zll_main_finishinstr1_in = arg0;
  assign zll_main_putaddrout1_in = {zll_main_finishinstr1_in[75:70], zll_main_finishinstr1_in[69:0]};
  ZLL_Main_putAddrOut1  inst (zll_main_putaddrout1_in[75:70], zll_main_putaddrout1_in[69:0], zll_main_putaddrout1_out);
  assign main_putweout_in = zll_main_putaddrout1_out;
  Main_putWeOut  instR1 (main_putweout_in[69:0], main_putweout_out);
  assign res = main_putweout_out;
endmodule

module Main_getOut (input logic [69:0] arg0,
  output logic [84:0] res);
  logic [139:0] zll_main_getout_in;
  logic [139:0] zll_main_getout1_in;
  logic [69:0] zll_main_outputs6_in;
  logic [69:0] zll_main_outputs2_in;
  logic [61:0] zll_main_outputs3_in;
  logic [53:0] zll_main_outputs4_in;
  logic [45:0] zll_main_outputs5_in;
  logic [37:0] zll_main_outputs_in;
  logic [31:0] zll_main_outputs7_in;
  assign zll_main_getout_in = {arg0, arg0};
  assign zll_main_getout1_in = zll_main_getout_in[139:0];
  assign zll_main_outputs6_in = zll_main_getout1_in[139:70];
  assign zll_main_outputs2_in = zll_main_outputs6_in[69:0];
  assign zll_main_outputs3_in = {zll_main_outputs2_in[61:54], zll_main_outputs2_in[53:46], zll_main_outputs2_in[45:38], zll_main_outputs2_in[37:32], zll_main_outputs2_in[31:15], zll_main_outputs2_in[14:0]};
  assign zll_main_outputs4_in = {zll_main_outputs3_in[53:46], zll_main_outputs3_in[45:38], zll_main_outputs3_in[37:32], zll_main_outputs3_in[31:15], zll_main_outputs3_in[14:0]};
  assign zll_main_outputs5_in = {zll_main_outputs4_in[45:38], zll_main_outputs4_in[37:32], zll_main_outputs4_in[31:15], zll_main_outputs4_in[14:0]};
  assign zll_main_outputs_in = {zll_main_outputs5_in[37:32], zll_main_outputs5_in[31:15], zll_main_outputs5_in[14:0]};
  assign zll_main_outputs7_in = {zll_main_outputs_in[31:15], zll_main_outputs_in[14:0]};
  assign res = {zll_main_outputs7_in[14:0], zll_main_getout1_in[69:0]};
endmodule

module ZLL_Main_r13 (input logic [7:0] arg0,
  input logic [7:0] arg1,
  input logic [7:0] arg2,
  input logic [5:0] arg3,
  input logic [16:0] arg4,
  input logic [14:0] arg5,
  output logic [7:0] res);
  logic [53:0] zll_main_r27_in;
  logic [7:0] zll_main_r27_out;
  assign zll_main_r27_in = {arg0, arg2, arg3, arg4, arg5};
  ZLL_Main_r27  inst (zll_main_r27_in[53:46], zll_main_r27_in[45:38], zll_main_r27_in[37:32], zll_main_r27_in[31:15], zll_main_r27_in[14:0], zll_main_r27_out);
  assign res = zll_main_r27_out;
endmodule

module ZLL_Main_putReg27 (input logic [7:0] arg0,
  input logic [1:0] arg1,
  input logic [9:0] arg2,
  input logic [69:0] arg3,
  output logic [69:0] res);
  logic [89:0] zll_main_putreg57_in;
  logic [89:0] zll_main_putreg25_in;
  logic [79:0] zll_main_putreg40_in;
  logic [79:0] zll_main_putreg18_in;
  logic [77:0] zll_main_putreg55_in;
  logic [77:0] zll_main_putreg16_in;
  logic [147:0] zll_main_putreg53_in;
  logic [147:0] zll_main_putreg48_in;
  logic [77:0] zll_main_putreg37_in;
  logic [77:0] zll_main_putreg13_in;
  logic [77:0] zll_main_putreg64_in;
  logic [77:0] zll_main_putreg35_in;
  logic [69:0] zll_main_putreg4_in;
  logic [79:0] zll_main_putreg36_in;
  logic [77:0] zll_main_putreg10_in;
  logic [77:0] zll_main_putreg33_in;
  logic [147:0] zll_main_putreg32_in;
  logic [147:0] zll_main_putreg43_in;
  logic [77:0] zll_main_putreg28_in;
  logic [77:0] zll_main_putreg67_in;
  logic [77:0] zll_main_putreg14_in;
  logic [69:0] zll_main_putreg20_in;
  logic [69:0] zll_main_putreg22_in;
  logic [79:0] zll_main_putreg52_in;
  logic [77:0] zll_main_putreg7_in;
  logic [77:0] zll_main_putreg58_in;
  logic [147:0] zll_main_putreg46_in;
  logic [147:0] zll_main_putreg51_in;
  logic [77:0] zll_main_putreg5_in;
  logic [77:0] zll_main_putreg42_in;
  logic [77:0] zll_main_putreg29_in;
  logic [69:0] zll_main_putreg62_in;
  logic [69:0] zll_main_putreg17_in;
  logic [69:0] zll_main_putreg24_in;
  logic [79:0] zll_main_putreg11_in;
  logic [77:0] zll_main_putreg61_in;
  logic [77:0] zll_main_putreg63_in;
  logic [147:0] zll_main_putreg21_in;
  logic [147:0] zll_main_putreg59_in;
  logic [77:0] zll_main_putreg2_in;
  logic [77:0] zll_main_putreg66_in;
  logic [69:0] zll_main_putreg47_in;
  logic [69:0] zll_main_putreg19_in;
  logic [69:0] zll_main_putreg49_in;
  logic [69:0] zll_main_putreg_in;
  assign zll_main_putreg57_in = {arg0, arg1, arg1, arg0, arg3};
  assign zll_main_putreg25_in = {zll_main_putreg57_in[89:82], zll_main_putreg57_in[81:80], zll_main_putreg57_in[81:80], zll_main_putreg57_in[89:82], zll_main_putreg57_in[69:0]};
  assign zll_main_putreg40_in = {zll_main_putreg25_in[81:80], zll_main_putreg25_in[89:82], zll_main_putreg25_in[69:0]};
  assign zll_main_putreg18_in = {zll_main_putreg40_in[69:0], zll_main_putreg40_in[79:70]};
  assign zll_main_putreg55_in = {zll_main_putreg18_in[79:10], zll_main_putreg18_in[7:0]};
  assign zll_main_putreg16_in = {zll_main_putreg55_in[7:0], zll_main_putreg55_in[77:8]};
  assign zll_main_putreg53_in = {zll_main_putreg16_in[77:70], zll_main_putreg16_in[69:0], zll_main_putreg16_in[69:0]};
  assign zll_main_putreg48_in = {zll_main_putreg53_in[147:140], zll_main_putreg53_in[139:0]};
  assign zll_main_putreg37_in = {zll_main_putreg48_in[147:140], zll_main_putreg48_in[139:70]};
  assign zll_main_putreg13_in = {zll_main_putreg37_in[77:70], zll_main_putreg37_in[69:0]};
  assign zll_main_putreg64_in = {zll_main_putreg13_in[61:54], zll_main_putreg13_in[77:70], zll_main_putreg13_in[69:62], zll_main_putreg13_in[53:46], zll_main_putreg13_in[45:38], zll_main_putreg13_in[37:32], zll_main_putreg13_in[31:15], zll_main_putreg13_in[14:0]};
  assign zll_main_putreg35_in = {zll_main_putreg64_in[53:46], zll_main_putreg64_in[77:70], zll_main_putreg64_in[69:62], zll_main_putreg64_in[61:54], zll_main_putreg64_in[45:38], zll_main_putreg64_in[37:32], zll_main_putreg64_in[31:15], zll_main_putreg64_in[14:0]};
  assign zll_main_putreg4_in = {zll_main_putreg35_in[77:70], zll_main_putreg35_in[69:62], zll_main_putreg35_in[61:54], zll_main_putreg35_in[53:46], zll_main_putreg35_in[37:32], zll_main_putreg35_in[31:15], zll_main_putreg35_in[14:0]};
  assign zll_main_putreg36_in = {zll_main_putreg25_in[69:0], zll_main_putreg25_in[79:70]};
  assign zll_main_putreg10_in = {zll_main_putreg36_in[79:10], zll_main_putreg36_in[7:0]};
  assign zll_main_putreg33_in = {zll_main_putreg10_in[7:0], zll_main_putreg10_in[77:8]};
  assign zll_main_putreg32_in = {zll_main_putreg33_in[77:70], zll_main_putreg33_in[69:0], zll_main_putreg33_in[69:0]};
  assign zll_main_putreg43_in = {zll_main_putreg32_in[147:140], zll_main_putreg32_in[139:0]};
  assign zll_main_putreg28_in = {zll_main_putreg43_in[147:140], zll_main_putreg43_in[139:70]};
  assign zll_main_putreg67_in = {zll_main_putreg28_in[77:70], zll_main_putreg28_in[69:0]};
  assign zll_main_putreg14_in = {zll_main_putreg67_in[69:62], zll_main_putreg67_in[77:70], zll_main_putreg67_in[61:54], zll_main_putreg67_in[53:46], zll_main_putreg67_in[45:38], zll_main_putreg67_in[37:32], zll_main_putreg67_in[31:15], zll_main_putreg67_in[14:0]};
  assign zll_main_putreg20_in = {zll_main_putreg14_in[77:70], zll_main_putreg14_in[69:62], zll_main_putreg14_in[61:54], zll_main_putreg14_in[45:38], zll_main_putreg14_in[37:32], zll_main_putreg14_in[31:15], zll_main_putreg14_in[14:0]};
  assign zll_main_putreg22_in = {zll_main_putreg20_in[69:62], zll_main_putreg20_in[45:38], zll_main_putreg20_in[61:54], zll_main_putreg20_in[53:46], zll_main_putreg20_in[37:32], zll_main_putreg20_in[31:15], zll_main_putreg20_in[14:0]};
  assign zll_main_putreg52_in = {zll_main_putreg57_in[69:0], zll_main_putreg57_in[79:70]};
  assign zll_main_putreg7_in = {zll_main_putreg52_in[79:10], zll_main_putreg52_in[7:0]};
  assign zll_main_putreg58_in = {zll_main_putreg7_in[7:0], zll_main_putreg7_in[77:8]};
  assign zll_main_putreg46_in = {zll_main_putreg58_in[77:70], zll_main_putreg58_in[69:0], zll_main_putreg58_in[69:0]};
  assign zll_main_putreg51_in = {zll_main_putreg46_in[147:140], zll_main_putreg46_in[139:0]};
  assign zll_main_putreg5_in = {zll_main_putreg51_in[147:140], zll_main_putreg51_in[139:70]};
  assign zll_main_putreg42_in = {zll_main_putreg5_in[77:70], zll_main_putreg5_in[69:0]};
  assign zll_main_putreg29_in = {zll_main_putreg42_in[69:62], zll_main_putreg42_in[77:70], zll_main_putreg42_in[61:54], zll_main_putreg42_in[53:46], zll_main_putreg42_in[45:38], zll_main_putreg42_in[37:32], zll_main_putreg42_in[31:15], zll_main_putreg42_in[14:0]};
  assign zll_main_putreg62_in = {zll_main_putreg29_in[77:70], zll_main_putreg29_in[69:62], zll_main_putreg29_in[53:46], zll_main_putreg29_in[45:38], zll_main_putreg29_in[37:32], zll_main_putreg29_in[31:15], zll_main_putreg29_in[14:0]};
  assign zll_main_putreg17_in = {zll_main_putreg62_in[69:62], zll_main_putreg62_in[61:54], zll_main_putreg62_in[45:38], zll_main_putreg62_in[53:46], zll_main_putreg62_in[37:32], zll_main_putreg62_in[31:15], zll_main_putreg62_in[14:0]};
  assign zll_main_putreg24_in = {zll_main_putreg17_in[69:62], zll_main_putreg17_in[37:32], zll_main_putreg17_in[61:54], zll_main_putreg17_in[53:46], zll_main_putreg17_in[45:38], zll_main_putreg17_in[31:15], zll_main_putreg17_in[14:0]};
  assign zll_main_putreg11_in = {arg3, arg2};
  assign zll_main_putreg61_in = {zll_main_putreg11_in[79:10], zll_main_putreg11_in[7:0]};
  assign zll_main_putreg63_in = {zll_main_putreg61_in[7:0], zll_main_putreg61_in[77:8]};
  assign zll_main_putreg21_in = {zll_main_putreg63_in[77:70], zll_main_putreg63_in[69:0], zll_main_putreg63_in[69:0]};
  assign zll_main_putreg59_in = {zll_main_putreg21_in[147:140], zll_main_putreg21_in[139:0]};
  assign zll_main_putreg2_in = {zll_main_putreg59_in[147:140], zll_main_putreg59_in[139:70]};
  assign zll_main_putreg66_in = {zll_main_putreg2_in[77:70], zll_main_putreg2_in[69:0]};
  assign zll_main_putreg47_in = {zll_main_putreg66_in[77:70], zll_main_putreg66_in[61:54], zll_main_putreg66_in[53:46], zll_main_putreg66_in[45:38], zll_main_putreg66_in[37:32], zll_main_putreg66_in[31:15], zll_main_putreg66_in[14:0]};
  assign zll_main_putreg19_in = {zll_main_putreg47_in[61:54], zll_main_putreg47_in[69:62], zll_main_putreg47_in[53:46], zll_main_putreg47_in[45:38], zll_main_putreg47_in[37:32], zll_main_putreg47_in[31:15], zll_main_putreg47_in[14:0]};
  assign zll_main_putreg49_in = {zll_main_putreg19_in[69:62], zll_main_putreg19_in[53:46], zll_main_putreg19_in[61:54], zll_main_putreg19_in[45:38], zll_main_putreg19_in[37:32], zll_main_putreg19_in[31:15], zll_main_putreg19_in[14:0]};
  assign zll_main_putreg_in = {zll_main_putreg49_in[69:62], zll_main_putreg49_in[61:54], zll_main_putreg49_in[37:32], zll_main_putreg49_in[53:46], zll_main_putreg49_in[45:38], zll_main_putreg49_in[31:15], zll_main_putreg49_in[14:0]};
  assign res = (zll_main_putreg11_in[9:8] == 2'h0) ? {zll_main_putreg_in[47:40], zll_main_putreg_in[69:62], zll_main_putreg_in[61:54], zll_main_putreg_in[39:32], zll_main_putreg_in[53:48], zll_main_putreg_in[31:15], zll_main_putreg_in[14:0]} : ((zll_main_putreg52_in[9:8] == 2'h1) ? {zll_main_putreg24_in[69:62], zll_main_putreg24_in[55:48], zll_main_putreg24_in[39:32], zll_main_putreg24_in[47:40], zll_main_putreg24_in[61:56], zll_main_putreg24_in[31:15], zll_main_putreg24_in[14:0]} : ((zll_main_putreg36_in[9:8] == 2'h2) ? {zll_main_putreg22_in[69:62], zll_main_putreg22_in[45:38], zll_main_putreg22_in[53:46], zll_main_putreg22_in[61:54], zll_main_putreg22_in[37:32], zll_main_putreg22_in[31:15], zll_main_putreg22_in[14:0]} : {zll_main_putreg4_in[45:38], zll_main_putreg4_in[61:54], zll_main_putreg4_in[69:62], zll_main_putreg4_in[53:46], zll_main_putreg4_in[37:32], zll_main_putreg4_in[31:15], zll_main_putreg4_in[14:0]}));
endmodule

module ZLL_Main_putOut5 (input logic [14:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [154:0] zll_main_putout14_in;
  logic [154:0] zll_main_putout10_in;
  logic [84:0] zll_main_putout1_in;
  logic [84:0] zll_main_putout12_in;
  logic [84:0] zll_main_putout11_in;
  logic [84:0] zll_main_putout4_in;
  logic [84:0] zll_main_putout9_in;
  logic [84:0] zll_main_putout7_in;
  assign zll_main_putout14_in = {arg0, arg1, arg1};
  assign zll_main_putout10_in = {zll_main_putout14_in[154:140], zll_main_putout14_in[139:0]};
  assign zll_main_putout1_in = {zll_main_putout10_in[154:140], zll_main_putout10_in[139:70]};
  assign zll_main_putout12_in = {zll_main_putout1_in[84:70], zll_main_putout1_in[69:0]};
  assign zll_main_putout11_in = {zll_main_putout12_in[53:46], zll_main_putout12_in[84:70], zll_main_putout12_in[69:62], zll_main_putout12_in[61:54], zll_main_putout12_in[45:38], zll_main_putout12_in[37:32], zll_main_putout12_in[31:15], zll_main_putout12_in[14:0]};
  assign zll_main_putout4_in = {zll_main_putout11_in[84:77], zll_main_putout11_in[45:38], zll_main_putout11_in[76:62], zll_main_putout11_in[61:54], zll_main_putout11_in[53:46], zll_main_putout11_in[37:32], zll_main_putout11_in[31:15], zll_main_putout11_in[14:0]};
  assign zll_main_putout9_in = {zll_main_putout4_in[84:77], zll_main_putout4_in[37:32], zll_main_putout4_in[76:69], zll_main_putout4_in[68:54], zll_main_putout4_in[53:46], zll_main_putout4_in[45:38], zll_main_putout4_in[31:15], zll_main_putout4_in[14:0]};
  assign zll_main_putout7_in = {zll_main_putout9_in[84:77], zll_main_putout9_in[76:71], zll_main_putout9_in[31:15], zll_main_putout9_in[70:63], zll_main_putout9_in[62:48], zll_main_putout9_in[47:40], zll_main_putout9_in[39:32], zll_main_putout9_in[14:0]};
  assign res = {zll_main_putout7_in[30:23], zll_main_putout7_in[22:15], zll_main_putout7_in[84:77], zll_main_putout7_in[53:46], zll_main_putout7_in[76:71], zll_main_putout7_in[70:54], zll_main_putout7_in[45:31]};
endmodule

module Main_putWeOut (input logic [69:0] arg0,
  output logic [69:0] res);
  logic [70:0] zll_main_putweout2_in;
  logic [69:0] zll_main_putweout2_out;
  assign zll_main_putweout2_in = {1'h0, arg0};
  ZLL_Main_putWeOut2  inst (zll_main_putweout2_in[70], zll_main_putweout2_in[69:0], zll_main_putweout2_out);
  assign res = zll_main_putweout2_out;
endmodule

module ZLL_Main_putAddrOut1 (input logic [5:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [69:0] main_getout_in;
  logic [84:0] main_getout_out;
  logic [90:0] zll_main_putaddrout10_in;
  logic [90:0] zll_main_putaddrout9_in;
  logic [20:0] zll_main_putaddrout3_in;
  logic [20:0] zll_main_putaddrout6_in;
  logic [84:0] zll_main_putout5_in;
  logic [69:0] zll_main_putout5_out;
  assign main_getout_in = arg1;
  Main_getOut  inst (main_getout_in[69:0], main_getout_out);
  assign zll_main_putaddrout10_in = {arg0, main_getout_out};
  assign zll_main_putaddrout9_in = {zll_main_putaddrout10_in[90:85], zll_main_putaddrout10_in[84:0]};
  assign zll_main_putaddrout3_in = {zll_main_putaddrout9_in[90:85], zll_main_putaddrout9_in[84:70]};
  assign zll_main_putaddrout6_in = {zll_main_putaddrout3_in[20:15], zll_main_putaddrout3_in[14:0]};
  assign zll_main_putout5_in = {{zll_main_putaddrout6_in[14], zll_main_putaddrout6_in[20:15], zll_main_putaddrout6_in[7:0]}, zll_main_putaddrout9_in[69:0]};
  ZLL_Main_putOut5  instR1 (zll_main_putout5_in[84:70], zll_main_putout5_in[69:0], zll_main_putout5_out);
  assign res = zll_main_putout5_out;
endmodule

module ZLL_Main_putWeOut2 (input logic [0:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [69:0] main_getout_in;
  logic [84:0] main_getout_out;
  logic [85:0] zll_main_putweout10_in;
  logic [85:0] zll_main_putweout3_in;
  logic [15:0] zll_main_putweout8_in;
  logic [15:0] zll_main_putweout_in;
  logic [84:0] zll_main_putout5_in;
  logic [69:0] zll_main_putout5_out;
  assign main_getout_in = arg1;
  Main_getOut  inst (main_getout_in[69:0], main_getout_out);
  assign zll_main_putweout10_in = {arg0, main_getout_out};
  assign zll_main_putweout3_in = {zll_main_putweout10_in[85], zll_main_putweout10_in[84:0]};
  assign zll_main_putweout8_in = {zll_main_putweout3_in[85], zll_main_putweout3_in[84:70]};
  assign zll_main_putweout_in = {zll_main_putweout8_in[15], zll_main_putweout8_in[14:0]};
  assign zll_main_putout5_in = {{zll_main_putweout_in[15], zll_main_putweout_in[13:8], zll_main_putweout_in[7:0]}, zll_main_putweout3_in[69:0]};
  ZLL_Main_putOut5  instR1 (zll_main_putout5_in[84:70], zll_main_putout5_in[69:0], zll_main_putout5_out);
  assign res = zll_main_putout5_out;
endmodule

module Main_incrPC (input logic [69:0] arg0,
  output logic [69:0] res);
  logic [69:0] main_getpc_in;
  logic [75:0] main_getpc_out;
  logic [75:0] zll_main_incrpc1_in;
  logic [75:0] zll_main_incrpc_in;
  logic [11:0] binop_in;
  logic [75:0] zll_main_putpc14_in;
  logic [69:0] zll_main_putpc14_out;
  assign main_getpc_in = arg0;
  Main_getPC  inst (main_getpc_in[69:0], main_getpc_out);
  assign zll_main_incrpc1_in = main_getpc_out;
  assign zll_main_incrpc_in = zll_main_incrpc1_in[75:0];
  assign binop_in = {zll_main_incrpc_in[75:70], 6'h1};
  assign zll_main_putpc14_in = {binop_in[11:6] + binop_in[5:0], zll_main_incrpc_in[69:0]};
  ZLL_Main_putPC14  instR1 (zll_main_putpc14_in[75:70], zll_main_putpc14_in[69:0], zll_main_putpc14_out);
  assign res = zll_main_putpc14_out;
endmodule

module ZLL_Main_getReg6 (input logic [1:0] arg0,
  input logic [1:0] arg1,
  input logic [69:0] arg2,
  output logic [77:0] res);
  logic [73:0] zll_main_getreg13_in;
  logic [73:0] zll_main_getreg3_in;
  logic [71:0] zll_main_getreg12_in;
  logic [71:0] zll_main_getreg_in;
  logic [69:0] zll_main_getreg21_in;
  logic [139:0] zll_main_getreg11_in;
  logic [139:0] zll_main_getreg14_in;
  logic [69:0] zll_main_r34_in;
  logic [69:0] zll_main_r33_in;
  logic [61:0] zll_main_r3_in;
  logic [53:0] zll_main_r37_in;
  logic [45:0] zll_main_r35_in;
  logic [7:0] zll_main_r35_out;
  logic [71:0] zll_main_getreg9_in;
  logic [69:0] zll_main_getreg4_in;
  logic [139:0] zll_main_getreg16_in;
  logic [139:0] zll_main_getreg20_in;
  logic [69:0] zll_main_r24_in;
  logic [69:0] zll_main_r22_in;
  logic [61:0] zll_main_r23_in;
  logic [53:0] zll_main_r27_in;
  logic [7:0] zll_main_r27_out;
  logic [71:0] zll_main_getreg7_in;
  logic [69:0] zll_main_getreg10_in;
  logic [139:0] zll_main_getreg2_in;
  logic [139:0] zll_main_getreg18_in;
  logic [69:0] zll_main_r15_in;
  logic [69:0] zll_main_r14_in;
  logic [61:0] zll_main_r13_in;
  logic [7:0] zll_main_r13_out;
  logic [71:0] zll_main_getreg1_in;
  logic [69:0] zll_main_getreg22_in;
  logic [139:0] zll_main_getreg17_in;
  logic [139:0] zll_main_getreg15_in;
  logic [69:0] zll_main_r0_in;
  logic [69:0] zll_main_r05_in;
  logic [61:0] zll_main_r13_inR1;
  logic [7:0] zll_main_r13_outR1;
  assign zll_main_getreg13_in = {arg0, arg0, arg2};
  assign zll_main_getreg3_in = {zll_main_getreg13_in[73:72], zll_main_getreg13_in[73:72], zll_main_getreg13_in[69:0]};
  assign zll_main_getreg12_in = {zll_main_getreg3_in[73:72], zll_main_getreg3_in[69:0]};
  assign zll_main_getreg_in = {zll_main_getreg12_in[69:0], zll_main_getreg12_in[71:70]};
  assign zll_main_getreg21_in = zll_main_getreg_in[71:2];
  assign zll_main_getreg11_in = {zll_main_getreg21_in[69:0], zll_main_getreg21_in[69:0]};
  assign zll_main_getreg14_in = zll_main_getreg11_in[139:0];
  assign zll_main_r34_in = zll_main_getreg14_in[139:70];
  assign zll_main_r33_in = zll_main_r34_in[69:0];
  assign zll_main_r3_in = {zll_main_r33_in[61:54], zll_main_r33_in[53:46], zll_main_r33_in[45:38], zll_main_r33_in[37:32], zll_main_r33_in[31:15], zll_main_r33_in[14:0]};
  assign zll_main_r37_in = {zll_main_r3_in[53:46], zll_main_r3_in[45:38], zll_main_r3_in[37:32], zll_main_r3_in[31:15], zll_main_r3_in[14:0]};
  assign zll_main_r35_in = {zll_main_r37_in[45:38], zll_main_r37_in[37:32], zll_main_r37_in[31:15], zll_main_r37_in[14:0]};
  ZLL_Main_r35  inst (zll_main_r35_in[45:38], zll_main_r35_in[37:32], zll_main_r35_in[31:15], zll_main_r35_in[14:0], zll_main_r35_out);
  assign zll_main_getreg9_in = {zll_main_getreg3_in[69:0], zll_main_getreg3_in[71:70]};
  assign zll_main_getreg4_in = zll_main_getreg9_in[71:2];
  assign zll_main_getreg16_in = {zll_main_getreg4_in[69:0], zll_main_getreg4_in[69:0]};
  assign zll_main_getreg20_in = zll_main_getreg16_in[139:0];
  assign zll_main_r24_in = zll_main_getreg20_in[139:70];
  assign zll_main_r22_in = zll_main_r24_in[69:0];
  assign zll_main_r23_in = {zll_main_r22_in[61:54], zll_main_r22_in[53:46], zll_main_r22_in[45:38], zll_main_r22_in[37:32], zll_main_r22_in[31:15], zll_main_r22_in[14:0]};
  assign zll_main_r27_in = {zll_main_r23_in[53:46], zll_main_r23_in[45:38], zll_main_r23_in[37:32], zll_main_r23_in[31:15], zll_main_r23_in[14:0]};
  ZLL_Main_r27  instR1 (zll_main_r27_in[53:46], zll_main_r27_in[45:38], zll_main_r27_in[37:32], zll_main_r27_in[31:15], zll_main_r27_in[14:0], zll_main_r27_out);
  assign zll_main_getreg7_in = {zll_main_getreg13_in[69:0], zll_main_getreg13_in[71:70]};
  assign zll_main_getreg10_in = zll_main_getreg7_in[71:2];
  assign zll_main_getreg2_in = {zll_main_getreg10_in[69:0], zll_main_getreg10_in[69:0]};
  assign zll_main_getreg18_in = zll_main_getreg2_in[139:0];
  assign zll_main_r15_in = zll_main_getreg18_in[139:70];
  assign zll_main_r14_in = zll_main_r15_in[69:0];
  assign zll_main_r13_in = {zll_main_r14_in[61:54], zll_main_r14_in[53:46], zll_main_r14_in[45:38], zll_main_r14_in[37:32], zll_main_r14_in[31:15], zll_main_r14_in[14:0]};
  ZLL_Main_r13  instR2 (zll_main_r13_in[61:54], zll_main_r13_in[53:46], zll_main_r13_in[45:38], zll_main_r13_in[37:32], zll_main_r13_in[31:15], zll_main_r13_in[14:0], zll_main_r13_out);
  assign zll_main_getreg1_in = {arg2, arg1};
  assign zll_main_getreg22_in = zll_main_getreg1_in[71:2];
  assign zll_main_getreg17_in = {zll_main_getreg22_in[69:0], zll_main_getreg22_in[69:0]};
  assign zll_main_getreg15_in = zll_main_getreg17_in[139:0];
  assign zll_main_r0_in = zll_main_getreg15_in[139:70];
  assign zll_main_r05_in = zll_main_r0_in[69:0];
  assign zll_main_r13_inR1 = {zll_main_r05_in[69:62], zll_main_r05_in[53:46], zll_main_r05_in[45:38], zll_main_r05_in[37:32], zll_main_r05_in[31:15], zll_main_r05_in[14:0]};
  ZLL_Main_r13  instR3 (zll_main_r13_inR1[61:54], zll_main_r13_inR1[53:46], zll_main_r13_inR1[45:38], zll_main_r13_inR1[37:32], zll_main_r13_inR1[31:15], zll_main_r13_inR1[14:0], zll_main_r13_outR1);
  assign res = (zll_main_getreg1_in[1:0] == 2'h0) ? {zll_main_r13_outR1, zll_main_getreg15_in[69:0]} : ((zll_main_getreg7_in[1:0] == 2'h1) ? {zll_main_r13_out, zll_main_getreg18_in[69:0]} : ((zll_main_getreg9_in[1:0] == 2'h2) ? {zll_main_r27_out, zll_main_getreg20_in[69:0]} : {zll_main_r35_out, zll_main_getreg14_in[69:0]}));
endmodule

module Main_getPC (input logic [69:0] arg0,
  output logic [75:0] res);
  logic [139:0] zll_main_getpc1_in;
  logic [139:0] zll_main_getpc_in;
  logic [69:0] zll_main_pc6_in;
  logic [69:0] zll_main_pc3_in;
  logic [61:0] zll_main_pc4_in;
  logic [53:0] zll_main_pc2_in;
  logic [45:0] zll_main_pc_in;
  logic [37:0] zll_main_pc5_in;
  logic [20:0] zll_main_pc1_in;
  assign zll_main_getpc1_in = {arg0, arg0};
  assign zll_main_getpc_in = zll_main_getpc1_in[139:0];
  assign zll_main_pc6_in = zll_main_getpc_in[139:70];
  assign zll_main_pc3_in = zll_main_pc6_in[69:0];
  assign zll_main_pc4_in = {zll_main_pc3_in[61:54], zll_main_pc3_in[53:46], zll_main_pc3_in[45:38], zll_main_pc3_in[37:32], zll_main_pc3_in[31:15], zll_main_pc3_in[14:0]};
  assign zll_main_pc2_in = {zll_main_pc4_in[53:46], zll_main_pc4_in[45:38], zll_main_pc4_in[37:32], zll_main_pc4_in[31:15], zll_main_pc4_in[14:0]};
  assign zll_main_pc_in = {zll_main_pc2_in[45:38], zll_main_pc2_in[37:32], zll_main_pc2_in[31:15], zll_main_pc2_in[14:0]};
  assign zll_main_pc5_in = {zll_main_pc_in[37:32], zll_main_pc_in[31:15], zll_main_pc_in[14:0]};
  assign zll_main_pc1_in = {zll_main_pc5_in[37:32], zll_main_pc5_in[14:0]};
  assign res = {zll_main_pc1_in[20:15], zll_main_getpc_in[69:0]};
endmodule