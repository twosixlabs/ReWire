module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [16:0] __in0,
  output logic [14:0] __out0);
  logic [90:0] zll_pure_dispatch8_in;
  logic [142:0] zll_pure_dispatch8_out;
  logic [90:0] zll_pure_dispatch_in;
  logic [86:0] zll_main_reset30_in;
  logic [86:0] main_putins_in;
  logic [69:0] main_putins_out;
  logic [69:0] zll_main_loop259_in;
  logic [142:0] zll_main_loop259_out;
  logic [142:0] zll_main_reset_in;
  logic [142:0] zll_main_reset43_in;
  logic [69:0] zll_main_reset42_in;
  logic [69:0] main_getpc_in;
  logic [75:0] main_getpc_out;
  logic [75:0] zll_main_loop247_in;
  logic [69:0] zll_main_loop247_out;
  logic [69:0] zll_main_loop259_inR1;
  logic [142:0] zll_main_loop259_outR1;
  logic [142:0] zll_main_reset5_in;
  logic [142:0] zll_main_reset10_in;
  logic [69:0] zll_main_reset36_in;
  logic [69:0] main_getout_in;
  logic [84:0] main_getout_out;
  logic [84:0] zll_main_loop260_in;
  logic [142:0] zll_main_loop260_out;
  logic [142:0] zll_main_reset35_in;
  logic [142:0] zll_main_reset13_in;
  logic [84:0] zll_main_reset26_in;
  logic [90:0] zll_pure_dispatch8_inR1;
  logic [142:0] zll_pure_dispatch8_outR1;
  logic [90:0] zll_pure_dispatch8_inR2;
  logic [142:0] zll_pure_dispatch8_outR2;
  logic [90:0] zll_pure_dispatch8_inR3;
  logic [142:0] zll_pure_dispatch8_outR3;
  logic [90:0] zll_pure_dispatch6_in;
  logic [86:0] zll_main_loop73_in;
  logic [86:0] main_putins_inR1;
  logic [69:0] main_putins_outR1;
  logic [69:0] zll_main_loop259_inR2;
  logic [142:0] zll_main_loop259_outR2;
  logic [142:0] zll_main_loop183_in;
  logic [142:0] zll_main_loop262_in;
  logic [69:0] zll_main_loop55_in;
  logic [69:0] main_incrpc_in;
  logic [69:0] main_incrpc_out;
  logic [69:0] zll_main_loop259_inR3;
  logic [142:0] zll_main_loop259_outR3;
  logic [142:0] zll_main_loop158_in;
  logic [142:0] zll_main_loop59_in;
  logic [69:0] zll_main_loop252_in;
  logic [69:0] main_getpc_inR1;
  logic [75:0] main_getpc_outR1;
  logic [75:0] zll_main_loop247_inR1;
  logic [69:0] zll_main_loop247_outR1;
  logic [69:0] zll_main_loop259_inR4;
  logic [142:0] zll_main_loop259_outR4;
  logic [142:0] zll_main_loop6_in;
  logic [142:0] zll_main_loop109_in;
  logic [69:0] zll_main_loop168_in;
  logic [69:0] main_getout_inR1;
  logic [84:0] main_getout_outR1;
  logic [84:0] zll_main_loop260_inR1;
  logic [142:0] zll_main_loop260_outR1;
  logic [142:0] zll_main_loop232_in;
  logic [142:0] zll_main_loop108_in;
  logic [84:0] zll_main_loop133_in;
  logic [90:0] zll_pure_dispatch8_inR4;
  logic [142:0] zll_pure_dispatch8_outR4;
  logic [90:0] zll_pure_dispatch1_in;
  logic [86:0] zll_main_loop136_in;
  logic [86:0] main_putins_inR2;
  logic [69:0] main_putins_outR2;
  logic [69:0] zll_main_loop259_inR5;
  logic [142:0] zll_main_loop259_outR5;
  logic [142:0] zll_main_loop66_in;
  logic [142:0] zll_main_loop38_in;
  logic [69:0] zll_main_loop112_in;
  logic [69:0] main_incrpc_inR1;
  logic [69:0] main_incrpc_outR1;
  logic [69:0] zll_main_loop259_inR6;
  logic [142:0] zll_main_loop259_outR6;
  logic [142:0] zll_main_loop179_in;
  logic [142:0] zll_main_loop261_in;
  logic [69:0] zll_main_loop43_in;
  logic [69:0] main_getpc_inR2;
  logic [75:0] main_getpc_outR2;
  logic [75:0] zll_main_loop247_inR2;
  logic [69:0] zll_main_loop247_outR2;
  logic [69:0] zll_main_loop259_inR7;
  logic [142:0] zll_main_loop259_outR7;
  logic [142:0] zll_main_loop240_in;
  logic [142:0] zll_main_loop145_in;
  logic [69:0] zll_main_loop42_in;
  logic [69:0] main_getout_inR2;
  logic [84:0] main_getout_outR2;
  logic [84:0] zll_main_loop260_inR2;
  logic [142:0] zll_main_loop260_outR2;
  logic [142:0] zll_main_loop130_in;
  logic [142:0] zll_main_loop142_in;
  logic [84:0] zll_main_loop116_in;
  logic [90:0] zll_pure_dispatch5_in;
  logic [86:0] zll_main_loop80_in;
  logic [86:0] main_putins_inR3;
  logic [69:0] main_putins_outR3;
  logic [69:0] zll_main_loop259_inR8;
  logic [142:0] zll_main_loop259_outR8;
  logic [142:0] zll_main_loop146_in;
  logic [142:0] zll_main_loop152_in;
  logic [69:0] zll_main_loop84_in;
  logic [69:0] main_getdatain_in;
  logic [69:0] main_getins_in;
  logic [86:0] main_getins_out;
  logic [86:0] zll_main_getdatain1_in;
  logic [86:0] zll_main_getdatain_in;
  logic [16:0] main_datain_in;
  logic [16:0] zll_main_datain_in;
  logic [77:0] zll_main_loop250_in;
  logic [77:0] main_putreg1_in;
  logic [69:0] main_putreg1_out;
  logic [69:0] zll_main_loop259_inR9;
  logic [142:0] zll_main_loop259_outR9;
  logic [142:0] zll_main_loop138_in;
  logic [142:0] zll_main_loop138_out;
  logic [0:0] __continue;
  logic [52:0] __padding;
  logic [3:0] __resumption_tag;
  logic [69:0] __st0;
  logic [3:0] __resumption_tag_next;
  logic [69:0] __st0_next;
  assign zll_pure_dispatch8_in = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch8  inst (zll_pure_dispatch8_in[90:74], zll_pure_dispatch8_in[69:0], zll_pure_dispatch8_out);
  assign zll_pure_dispatch_in = {__in0, {__resumption_tag, __st0}};
  assign zll_main_reset30_in = {zll_pure_dispatch_in[90:74], zll_pure_dispatch_in[69:0]};
  assign main_putins_in = {zll_main_reset30_in[86:70], zll_main_reset30_in[69:0]};
  Main_putIns  instR1 (main_putins_in[86:70], main_putins_in[69:0], main_putins_out);
  assign zll_main_loop259_in = main_putins_out;
  ZLL_Main_loop259  instR2 (zll_main_loop259_in[69:0], zll_main_loop259_out);
  assign zll_main_reset_in = zll_main_loop259_out;
  assign zll_main_reset43_in = zll_main_reset_in[142:0];
  assign zll_main_reset42_in = zll_main_reset43_in[69:0];
  assign main_getpc_in = zll_main_reset42_in[69:0];
  Main_getPC  instR3 (main_getpc_in[69:0], main_getpc_out);
  assign zll_main_loop247_in = main_getpc_out;
  ZLL_Main_loop247  instR4 (zll_main_loop247_in[75:0], zll_main_loop247_out);
  assign zll_main_loop259_inR1 = zll_main_loop247_out;
  ZLL_Main_loop259  instR5 (zll_main_loop259_inR1[69:0], zll_main_loop259_outR1);
  assign zll_main_reset5_in = zll_main_loop259_outR1;
  assign zll_main_reset10_in = zll_main_reset5_in[142:0];
  assign zll_main_reset36_in = zll_main_reset10_in[69:0];
  assign main_getout_in = zll_main_reset36_in[69:0];
  Main_getOut  instR6 (main_getout_in[69:0], main_getout_out);
  assign zll_main_loop260_in = main_getout_out;
  ZLL_Main_loop260  instR7 (zll_main_loop260_in[84:0], zll_main_loop260_out);
  assign zll_main_reset35_in = zll_main_loop260_out;
  assign zll_main_reset13_in = zll_main_reset35_in[142:0];
  assign zll_main_reset26_in = {zll_main_reset13_in[84:70], zll_main_reset13_in[69:0]};
  assign zll_pure_dispatch8_inR1 = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch8  instR8 (zll_pure_dispatch8_inR1[90:74], zll_pure_dispatch8_inR1[69:0], zll_pure_dispatch8_outR1);
  assign zll_pure_dispatch8_inR2 = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch8  instR9 (zll_pure_dispatch8_inR2[90:74], zll_pure_dispatch8_inR2[69:0], zll_pure_dispatch8_outR2);
  assign zll_pure_dispatch8_inR3 = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch8  instR10 (zll_pure_dispatch8_inR3[90:74], zll_pure_dispatch8_inR3[69:0], zll_pure_dispatch8_outR3);
  assign zll_pure_dispatch6_in = {__in0, {__resumption_tag, __st0}};
  assign zll_main_loop73_in = {zll_pure_dispatch6_in[90:74], zll_pure_dispatch6_in[69:0]};
  assign main_putins_inR1 = {zll_main_loop73_in[86:70], zll_main_loop73_in[69:0]};
  Main_putIns  instR11 (main_putins_inR1[86:70], main_putins_inR1[69:0], main_putins_outR1);
  assign zll_main_loop259_inR2 = main_putins_outR1;
  ZLL_Main_loop259  instR12 (zll_main_loop259_inR2[69:0], zll_main_loop259_outR2);
  assign zll_main_loop183_in = zll_main_loop259_outR2;
  assign zll_main_loop262_in = zll_main_loop183_in[142:0];
  assign zll_main_loop55_in = zll_main_loop262_in[69:0];
  assign main_incrpc_in = zll_main_loop55_in[69:0];
  Main_incrPC  instR13 (main_incrpc_in[69:0], main_incrpc_out);
  assign zll_main_loop259_inR3 = main_incrpc_out;
  ZLL_Main_loop259  instR14 (zll_main_loop259_inR3[69:0], zll_main_loop259_outR3);
  assign zll_main_loop158_in = zll_main_loop259_outR3;
  assign zll_main_loop59_in = zll_main_loop158_in[142:0];
  assign zll_main_loop252_in = zll_main_loop59_in[69:0];
  assign main_getpc_inR1 = zll_main_loop252_in[69:0];
  Main_getPC  instR15 (main_getpc_inR1[69:0], main_getpc_outR1);
  assign zll_main_loop247_inR1 = main_getpc_outR1;
  ZLL_Main_loop247  instR16 (zll_main_loop247_inR1[75:0], zll_main_loop247_outR1);
  assign zll_main_loop259_inR4 = zll_main_loop247_outR1;
  ZLL_Main_loop259  instR17 (zll_main_loop259_inR4[69:0], zll_main_loop259_outR4);
  assign zll_main_loop6_in = zll_main_loop259_outR4;
  assign zll_main_loop109_in = zll_main_loop6_in[142:0];
  assign zll_main_loop168_in = zll_main_loop109_in[69:0];
  assign main_getout_inR1 = zll_main_loop168_in[69:0];
  Main_getOut  instR18 (main_getout_inR1[69:0], main_getout_outR1);
  assign zll_main_loop260_inR1 = main_getout_outR1;
  ZLL_Main_loop260  instR19 (zll_main_loop260_inR1[84:0], zll_main_loop260_outR1);
  assign zll_main_loop232_in = zll_main_loop260_outR1;
  assign zll_main_loop108_in = zll_main_loop232_in[142:0];
  assign zll_main_loop133_in = {zll_main_loop108_in[84:70], zll_main_loop108_in[69:0]};
  assign zll_pure_dispatch8_inR4 = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch8  instR20 (zll_pure_dispatch8_inR4[90:74], zll_pure_dispatch8_inR4[69:0], zll_pure_dispatch8_outR4);
  assign zll_pure_dispatch1_in = {__in0, {__resumption_tag, __st0}};
  assign zll_main_loop136_in = {zll_pure_dispatch1_in[90:74], zll_pure_dispatch1_in[69:0]};
  assign main_putins_inR2 = {zll_main_loop136_in[86:70], zll_main_loop136_in[69:0]};
  Main_putIns  instR21 (main_putins_inR2[86:70], main_putins_inR2[69:0], main_putins_outR2);
  assign zll_main_loop259_inR5 = main_putins_outR2;
  ZLL_Main_loop259  instR22 (zll_main_loop259_inR5[69:0], zll_main_loop259_outR5);
  assign zll_main_loop66_in = zll_main_loop259_outR5;
  assign zll_main_loop38_in = zll_main_loop66_in[142:0];
  assign zll_main_loop112_in = zll_main_loop38_in[69:0];
  assign main_incrpc_inR1 = zll_main_loop112_in[69:0];
  Main_incrPC  instR23 (main_incrpc_inR1[69:0], main_incrpc_outR1);
  assign zll_main_loop259_inR6 = main_incrpc_outR1;
  ZLL_Main_loop259  instR24 (zll_main_loop259_inR6[69:0], zll_main_loop259_outR6);
  assign zll_main_loop179_in = zll_main_loop259_outR6;
  assign zll_main_loop261_in = zll_main_loop179_in[142:0];
  assign zll_main_loop43_in = zll_main_loop261_in[69:0];
  assign main_getpc_inR2 = zll_main_loop43_in[69:0];
  Main_getPC  instR25 (main_getpc_inR2[69:0], main_getpc_outR2);
  assign zll_main_loop247_inR2 = main_getpc_outR2;
  ZLL_Main_loop247  instR26 (zll_main_loop247_inR2[75:0], zll_main_loop247_outR2);
  assign zll_main_loop259_inR7 = zll_main_loop247_outR2;
  ZLL_Main_loop259  instR27 (zll_main_loop259_inR7[69:0], zll_main_loop259_outR7);
  assign zll_main_loop240_in = zll_main_loop259_outR7;
  assign zll_main_loop145_in = zll_main_loop240_in[142:0];
  assign zll_main_loop42_in = zll_main_loop145_in[69:0];
  assign main_getout_inR2 = zll_main_loop42_in[69:0];
  Main_getOut  instR28 (main_getout_inR2[69:0], main_getout_outR2);
  assign zll_main_loop260_inR2 = main_getout_outR2;
  ZLL_Main_loop260  instR29 (zll_main_loop260_inR2[84:0], zll_main_loop260_outR2);
  assign zll_main_loop130_in = zll_main_loop260_outR2;
  assign zll_main_loop142_in = zll_main_loop130_in[142:0];
  assign zll_main_loop116_in = {zll_main_loop142_in[84:70], zll_main_loop142_in[69:0]};
  assign zll_pure_dispatch5_in = {__in0, {__resumption_tag, __st0}};
  assign zll_main_loop80_in = {zll_pure_dispatch5_in[90:74], zll_pure_dispatch5_in[69:0]};
  assign main_putins_inR3 = {zll_main_loop80_in[86:70], zll_main_loop80_in[69:0]};
  Main_putIns  instR30 (main_putins_inR3[86:70], main_putins_inR3[69:0], main_putins_outR3);
  assign zll_main_loop259_inR8 = main_putins_outR3;
  ZLL_Main_loop259  instR31 (zll_main_loop259_inR8[69:0], zll_main_loop259_outR8);
  assign zll_main_loop146_in = zll_main_loop259_outR8;
  assign zll_main_loop152_in = zll_main_loop146_in[142:0];
  assign zll_main_loop84_in = zll_main_loop152_in[69:0];
  assign main_getdatain_in = zll_main_loop84_in[69:0];
  assign main_getins_in = main_getdatain_in[69:0];
  Main_getIns  instR32 (main_getins_in[69:0], main_getins_out);
  assign zll_main_getdatain1_in = main_getins_out;
  assign zll_main_getdatain_in = zll_main_getdatain1_in[86:0];
  assign main_datain_in = zll_main_getdatain_in[86:70];
  assign zll_main_datain_in = main_datain_in[16:0];
  assign zll_main_loop250_in = {zll_main_datain_in[7:0], zll_main_getdatain_in[69:0]};
  assign main_putreg1_in = zll_main_loop250_in[77:0];
  Main_putReg1  instR33 (main_putreg1_in[77:70], main_putreg1_in[69:0], main_putreg1_out);
  assign zll_main_loop259_inR9 = main_putreg1_out;
  ZLL_Main_loop259  instR34 (zll_main_loop259_inR9[69:0], zll_main_loop259_outR9);
  assign zll_main_loop138_in = zll_main_loop259_outR9;
  ZLL_Main_loop138  instR35 (zll_main_loop138_in[142:0], zll_main_loop138_out);
  assign {__continue, __padding, __out0, __resumption_tag_next, __st0_next} = (zll_pure_dispatch5_in[73:70] == 4'h1) ? zll_main_loop138_out : ((zll_pure_dispatch1_in[73:70] == 4'h2) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop116_in[84:70], 4'h1, zll_main_loop116_in[69:0]} : ((zll_pure_dispatch8_inR4[73:70] == 4'h3) ? zll_pure_dispatch8_outR4 : ((zll_pure_dispatch6_in[73:70] == 4'h4) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop133_in[84:70], 4'h3, zll_main_loop133_in[69:0]} : ((zll_pure_dispatch8_inR3[73:70] == 4'h5) ? zll_pure_dispatch8_outR3 : ((zll_pure_dispatch8_inR2[73:70] == 4'h6) ? zll_pure_dispatch8_outR2 : ((zll_pure_dispatch8_inR1[73:70] == 4'h7) ? zll_pure_dispatch8_outR1 : ((zll_pure_dispatch_in[73:70] == 4'h8) ? {{1'h1, {6'h35{1'h0}}}, zll_main_reset26_in[84:70], 4'h7, zll_main_reset26_in[69:0]} : zll_pure_dispatch8_out)))))));
  initial {__resumption_tag, __st0} <= {1'h1, {7'h49{1'h0}}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      {__resumption_tag, __st0} <= {1'h1, {7'h49{1'h0}}};
    end else begin
      {__resumption_tag, __st0} <= {__resumption_tag_next, __st0_next};
    end
  end
endmodule

module ZLL_Main_loop260 (input logic [84:0] arg0,
  output logic [142:0] res);
  logic [84:0] zll_main_loop244_in;
  assign zll_main_loop244_in = arg0;
  assign res = {{2'h1, {6'h38{1'h0}}}, zll_main_loop244_in[84:70], zll_main_loop244_in[69:0]};
endmodule

module ZLL_Main_loop259 (input logic [69:0] arg0,
  output logic [142:0] res);
  assign res = {{7'h49{1'h0}}, arg0};
endmodule

module ZLL_Pure_dispatch8 (input logic [16:0] arg0,
  input logic [69:0] arg1,
  output logic [142:0] res);
  logic [86:0] zll_main_loop249_in;
  logic [86:0] main_putins_in;
  logic [69:0] main_putins_out;
  logic [69:0] zll_main_loop259_in;
  logic [142:0] zll_main_loop259_out;
  logic [142:0] zll_main_loop138_in;
  logic [142:0] zll_main_loop138_out;
  assign zll_main_loop249_in = {arg0, arg1};
  assign main_putins_in = {zll_main_loop249_in[86:70], zll_main_loop249_in[69:0]};
  Main_putIns  inst (main_putins_in[86:70], main_putins_in[69:0], main_putins_out);
  assign zll_main_loop259_in = main_putins_out;
  ZLL_Main_loop259  instR1 (zll_main_loop259_in[69:0], zll_main_loop259_out);
  assign zll_main_loop138_in = zll_main_loop259_out;
  ZLL_Main_loop138  instR2 (zll_main_loop138_in[142:0], zll_main_loop138_out);
  assign res = zll_main_loop138_out;
endmodule

module ZLL_Main_loop247 (input logic [75:0] arg0,
  output logic [69:0] res);
  logic [75:0] zll_main_loop217_in;
  logic [75:0] main_putaddrout_in;
  logic [69:0] main_putaddrout_out;
  logic [69:0] main_putweout1_in;
  logic [69:0] main_putweout1_out;
  assign zll_main_loop217_in = arg0;
  assign main_putaddrout_in = {zll_main_loop217_in[75:70], zll_main_loop217_in[69:0]};
  Main_putAddrOut  inst (main_putaddrout_in[75:70], main_putaddrout_in[69:0], main_putaddrout_out);
  assign main_putweout1_in = main_putaddrout_out;
  Main_putWeOut1  instR1 (main_putweout1_in[69:0], main_putweout1_out);
  assign res = main_putweout1_out;
endmodule

module Main_putPC1 (input logic [5:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [145:0] zll_main_putpc10_in;
  logic [145:0] zll_main_putpc7_in;
  logic [75:0] zll_main_putpc3_in;
  logic [75:0] zll_main_putpc9_in;
  logic [75:0] zll_main_putpc8_in;
  logic [75:0] zll_main_putpc4_in;
  logic [75:0] zll_main_putpc12_in;
  assign zll_main_putpc10_in = {arg0, arg1, arg1};
  assign zll_main_putpc7_in = {zll_main_putpc10_in[145:140], zll_main_putpc10_in[139:0]};
  assign zll_main_putpc3_in = {zll_main_putpc7_in[145:140], zll_main_putpc7_in[139:70]};
  assign zll_main_putpc9_in = {zll_main_putpc3_in[69:62], zll_main_putpc3_in[75:70], zll_main_putpc3_in[61:54], zll_main_putpc3_in[53:46], zll_main_putpc3_in[45:38], zll_main_putpc3_in[37:32], zll_main_putpc3_in[31:15], zll_main_putpc3_in[14:0]};
  assign zll_main_putpc8_in = {zll_main_putpc9_in[75:68], zll_main_putpc9_in[61:54], zll_main_putpc9_in[67:62], zll_main_putpc9_in[53:46], zll_main_putpc9_in[45:38], zll_main_putpc9_in[37:32], zll_main_putpc9_in[31:15], zll_main_putpc9_in[14:0]};
  assign zll_main_putpc4_in = {zll_main_putpc8_in[75:68], zll_main_putpc8_in[53:46], zll_main_putpc8_in[67:60], zll_main_putpc8_in[59:54], zll_main_putpc8_in[45:38], zll_main_putpc8_in[37:32], zll_main_putpc8_in[31:15], zll_main_putpc8_in[14:0]};
  assign zll_main_putpc12_in = {zll_main_putpc4_in[75:68], zll_main_putpc4_in[45:38], zll_main_putpc4_in[67:60], zll_main_putpc4_in[59:52], zll_main_putpc4_in[51:46], zll_main_putpc4_in[37:32], zll_main_putpc4_in[31:15], zll_main_putpc4_in[14:0]};
  assign res = {zll_main_putpc12_in[75:68], zll_main_putpc12_in[51:44], zll_main_putpc12_in[59:52], zll_main_putpc12_in[67:60], zll_main_putpc12_in[43:38], zll_main_putpc12_in[31:15], zll_main_putpc12_in[14:0]};
endmodule

module Main_putIns (input logic [16:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [156:0] zll_main_putins9_in;
  logic [156:0] zll_main_putins5_in;
  logic [86:0] zll_main_putins10_in;
  logic [86:0] zll_main_putins1_in;
  logic [86:0] zll_main_putins4_in;
  logic [86:0] zll_main_putins3_in;
  assign zll_main_putins9_in = {arg0, arg1, arg1};
  assign zll_main_putins5_in = {zll_main_putins9_in[156:140], zll_main_putins9_in[139:0]};
  assign zll_main_putins10_in = {zll_main_putins5_in[156:140], zll_main_putins5_in[139:70]};
  assign zll_main_putins1_in = {zll_main_putins10_in[61:54], zll_main_putins10_in[86:70], zll_main_putins10_in[69:62], zll_main_putins10_in[53:46], zll_main_putins10_in[45:38], zll_main_putins10_in[37:32], zll_main_putins10_in[31:15], zll_main_putins10_in[14:0]};
  assign zll_main_putins4_in = {zll_main_putins1_in[86:79], zll_main_putins1_in[53:46], zll_main_putins1_in[78:62], zll_main_putins1_in[61:54], zll_main_putins1_in[45:38], zll_main_putins1_in[37:32], zll_main_putins1_in[31:15], zll_main_putins1_in[14:0]};
  assign zll_main_putins3_in = {zll_main_putins4_in[86:79], zll_main_putins4_in[78:71], zll_main_putins4_in[37:32], zll_main_putins4_in[70:54], zll_main_putins4_in[53:46], zll_main_putins4_in[45:38], zll_main_putins4_in[31:15], zll_main_putins4_in[14:0]};
  assign res = {zll_main_putins3_in[47:40], zll_main_putins3_in[86:79], zll_main_putins3_in[78:71], zll_main_putins3_in[39:32], zll_main_putins3_in[70:65], zll_main_putins3_in[64:48], zll_main_putins3_in[14:0]};
endmodule

module ZLL_Main_r06 (input logic [7:0] arg0,
  input logic [7:0] arg1,
  input logic [7:0] arg2,
  input logic [5:0] arg3,
  input logic [16:0] arg4,
  input logic [14:0] arg5,
  output logic [7:0] res);
  logic [53:0] zll_main_r14_in;
  logic [7:0] zll_main_r14_out;
  assign zll_main_r14_in = {arg0, arg2, arg3, arg4, arg5};
  ZLL_Main_r14  inst (zll_main_r14_in[53:46], zll_main_r14_in[45:38], zll_main_r14_in[37:32], zll_main_r14_in[31:15], zll_main_r14_in[14:0], zll_main_r14_out);
  assign res = zll_main_r14_out;
endmodule

module ZLL_Main_r14 (input logic [7:0] arg0,
  input logic [7:0] arg1,
  input logic [5:0] arg2,
  input logic [16:0] arg3,
  input logic [14:0] arg4,
  output logic [7:0] res);
  logic [45:0] zll_main_r26_in;
  logic [7:0] zll_main_r26_out;
  assign zll_main_r26_in = {arg0, arg2, arg3, arg4};
  ZLL_Main_r26  inst (zll_main_r26_in[45:38], zll_main_r26_in[37:32], zll_main_r26_in[31:15], zll_main_r26_in[14:0], zll_main_r26_out);
  assign res = zll_main_r26_out;
endmodule

module Main_putWeOut1 (input logic [69:0] arg0,
  output logic [69:0] res);
  logic [69:0] main_getout_in;
  logic [84:0] main_getout_out;
  logic [84:0] zll_main_putweout6_in;
  logic [84:0] zll_main_putweout4_in;
  logic [14:0] zll_main_putweout7_in;
  logic [84:0] main_putout_in;
  logic [69:0] main_putout_out;
  assign main_getout_in = arg0;
  Main_getOut  inst (main_getout_in[69:0], main_getout_out);
  assign zll_main_putweout6_in = main_getout_out;
  assign zll_main_putweout4_in = zll_main_putweout6_in[84:0];
  assign zll_main_putweout7_in = zll_main_putweout4_in[84:70];
  assign main_putout_in = {{1'h0, zll_main_putweout7_in[13:8], zll_main_putweout7_in[7:0]}, zll_main_putweout4_in[69:0]};
  Main_putOut  instR1 (main_putout_in[84:70], main_putout_in[69:0], main_putout_out);
  assign res = main_putout_out;
endmodule

module ZLL_Main_r26 (input logic [7:0] arg0,
  input logic [5:0] arg1,
  input logic [16:0] arg2,
  input logic [14:0] arg3,
  output logic [7:0] res);
  logic [39:0] zll_main_r16_in;
  logic [22:0] zll_main_r15_in;
  assign zll_main_r16_in = {arg0, arg2, arg3};
  assign zll_main_r15_in = {zll_main_r16_in[39:32], zll_main_r16_in[14:0]};
  assign res = zll_main_r15_in[22:15];
endmodule

module Main_getReg1 (input logic [1:0] arg0,
  input logic [69:0] arg1,
  output logic [77:0] res);
  logic [71:0] zll_main_getreg18_in;
  logic [69:0] zll_main_getreg10_in;
  logic [139:0] zll_main_getreg16_in;
  logic [139:0] zll_main_getreg5_in;
  logic [69:0] main_r3_in;
  logic [69:0] zll_main_r33_in;
  logic [61:0] zll_main_r32_in;
  logic [53:0] zll_main_r35_in;
  logic [45:0] zll_main_r26_in;
  logic [7:0] zll_main_r26_out;
  logic [71:0] zll_main_getreg4_in;
  logic [69:0] zll_main_getreg7_in;
  logic [139:0] zll_main_getreg1_in;
  logic [139:0] zll_main_getreg20_in;
  logic [69:0] main_r2_in;
  logic [69:0] zll_main_r23_in;
  logic [61:0] zll_main_r22_in;
  logic [53:0] zll_main_r14_in;
  logic [7:0] zll_main_r14_out;
  logic [71:0] zll_main_getreg9_in;
  logic [69:0] zll_main_getreg6_in;
  logic [139:0] zll_main_getreg_in;
  logic [139:0] zll_main_getreg15_in;
  logic [69:0] main_r1_in;
  logic [69:0] zll_main_r11_in;
  logic [61:0] zll_main_r06_in;
  logic [7:0] zll_main_r06_out;
  logic [71:0] zll_main_getreg21_in;
  logic [69:0] zll_main_getreg13_in;
  logic [77:0] zll_main_getreg13_out;
  assign zll_main_getreg18_in = {arg1, arg0};
  assign zll_main_getreg10_in = zll_main_getreg18_in[71:2];
  assign zll_main_getreg16_in = {zll_main_getreg10_in[69:0], zll_main_getreg10_in[69:0]};
  assign zll_main_getreg5_in = zll_main_getreg16_in[139:0];
  assign main_r3_in = zll_main_getreg5_in[139:70];
  assign zll_main_r33_in = main_r3_in[69:0];
  assign zll_main_r32_in = {zll_main_r33_in[61:54], zll_main_r33_in[53:46], zll_main_r33_in[45:38], zll_main_r33_in[37:32], zll_main_r33_in[31:15], zll_main_r33_in[14:0]};
  assign zll_main_r35_in = {zll_main_r32_in[53:46], zll_main_r32_in[45:38], zll_main_r32_in[37:32], zll_main_r32_in[31:15], zll_main_r32_in[14:0]};
  assign zll_main_r26_in = {zll_main_r35_in[45:38], zll_main_r35_in[37:32], zll_main_r35_in[31:15], zll_main_r35_in[14:0]};
  ZLL_Main_r26  inst (zll_main_r26_in[45:38], zll_main_r26_in[37:32], zll_main_r26_in[31:15], zll_main_r26_in[14:0], zll_main_r26_out);
  assign zll_main_getreg4_in = {arg1, arg0};
  assign zll_main_getreg7_in = zll_main_getreg4_in[71:2];
  assign zll_main_getreg1_in = {zll_main_getreg7_in[69:0], zll_main_getreg7_in[69:0]};
  assign zll_main_getreg20_in = zll_main_getreg1_in[139:0];
  assign main_r2_in = zll_main_getreg20_in[139:70];
  assign zll_main_r23_in = main_r2_in[69:0];
  assign zll_main_r22_in = {zll_main_r23_in[61:54], zll_main_r23_in[53:46], zll_main_r23_in[45:38], zll_main_r23_in[37:32], zll_main_r23_in[31:15], zll_main_r23_in[14:0]};
  assign zll_main_r14_in = {zll_main_r22_in[53:46], zll_main_r22_in[45:38], zll_main_r22_in[37:32], zll_main_r22_in[31:15], zll_main_r22_in[14:0]};
  ZLL_Main_r14  instR1 (zll_main_r14_in[53:46], zll_main_r14_in[45:38], zll_main_r14_in[37:32], zll_main_r14_in[31:15], zll_main_r14_in[14:0], zll_main_r14_out);
  assign zll_main_getreg9_in = {arg1, arg0};
  assign zll_main_getreg6_in = zll_main_getreg9_in[71:2];
  assign zll_main_getreg_in = {zll_main_getreg6_in[69:0], zll_main_getreg6_in[69:0]};
  assign zll_main_getreg15_in = zll_main_getreg_in[139:0];
  assign main_r1_in = zll_main_getreg15_in[139:70];
  assign zll_main_r11_in = main_r1_in[69:0];
  assign zll_main_r06_in = {zll_main_r11_in[61:54], zll_main_r11_in[53:46], zll_main_r11_in[45:38], zll_main_r11_in[37:32], zll_main_r11_in[31:15], zll_main_r11_in[14:0]};
  ZLL_Main_r06  instR2 (zll_main_r06_in[61:54], zll_main_r06_in[53:46], zll_main_r06_in[45:38], zll_main_r06_in[37:32], zll_main_r06_in[31:15], zll_main_r06_in[14:0], zll_main_r06_out);
  assign zll_main_getreg21_in = {arg1, arg0};
  assign zll_main_getreg13_in = zll_main_getreg21_in[71:2];
  ZLL_Main_getReg13  instR3 (zll_main_getreg13_in[69:0], zll_main_getreg13_out);
  assign res = (zll_main_getreg21_in[1:0] == 2'h0) ? zll_main_getreg13_out : ((zll_main_getreg9_in[1:0] == 2'h1) ? {zll_main_r06_out, zll_main_getreg15_in[69:0]} : ((zll_main_getreg4_in[1:0] == 2'h2) ? {zll_main_r14_out, zll_main_getreg20_in[69:0]} : {zll_main_r26_out, zll_main_getreg5_in[69:0]}));
endmodule

module Main_putReg1 (input logic [7:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [147:0] zll_main_putreg27_in;
  logic [147:0] zll_main_putreg36_in;
  logic [77:0] zll_main_putreg25_in;
  assign zll_main_putreg27_in = {arg0, arg1, arg1};
  assign zll_main_putreg36_in = {zll_main_putreg27_in[147:140], zll_main_putreg27_in[139:0]};
  assign zll_main_putreg25_in = {zll_main_putreg36_in[147:140], zll_main_putreg36_in[139:70]};
  assign res = {zll_main_putreg25_in[77:70], zll_main_putreg25_in[61:54], zll_main_putreg25_in[53:46], zll_main_putreg25_in[45:38], zll_main_putreg25_in[37:32], zll_main_putreg25_in[31:15], zll_main_putreg25_in[14:0]};
endmodule

module ZLL_Main_getReg13 (input logic [69:0] arg0,
  output logic [77:0] res);
  logic [139:0] zll_main_getreg19_in;
  logic [139:0] zll_main_getreg22_in;
  logic [69:0] main_r0_in;
  logic [69:0] zll_main_r03_in;
  logic [61:0] zll_main_r06_in;
  logic [7:0] zll_main_r06_out;
  assign zll_main_getreg19_in = {arg0, arg0};
  assign zll_main_getreg22_in = zll_main_getreg19_in[139:0];
  assign main_r0_in = zll_main_getreg22_in[139:70];
  assign zll_main_r03_in = main_r0_in[69:0];
  assign zll_main_r06_in = {zll_main_r03_in[69:62], zll_main_r03_in[53:46], zll_main_r03_in[45:38], zll_main_r03_in[37:32], zll_main_r03_in[31:15], zll_main_r03_in[14:0]};
  ZLL_Main_r06  inst (zll_main_r06_in[61:54], zll_main_r06_in[53:46], zll_main_r06_in[45:38], zll_main_r06_in[37:32], zll_main_r06_in[31:15], zll_main_r06_in[14:0], zll_main_r06_out);
  assign res = {zll_main_r06_out, zll_main_getreg22_in[69:0]};
endmodule

module Main_getIns (input logic [69:0] arg0,
  output logic [86:0] res);
  logic [139:0] zll_main_getins2_in;
  logic [139:0] zll_main_getins_in;
  logic [69:0] main_inputs_in;
  logic [69:0] zll_main_inputs_in;
  logic [61:0] zll_main_inputs2_in;
  logic [53:0] zll_main_inputs6_in;
  logic [45:0] zll_main_inputs3_in;
  logic [37:0] zll_main_inputs1_in;
  logic [31:0] zll_main_inputs4_in;
  assign zll_main_getins2_in = {arg0, arg0};
  assign zll_main_getins_in = zll_main_getins2_in[139:0];
  assign main_inputs_in = zll_main_getins_in[139:70];
  assign zll_main_inputs_in = main_inputs_in[69:0];
  assign zll_main_inputs2_in = {zll_main_inputs_in[61:54], zll_main_inputs_in[53:46], zll_main_inputs_in[45:38], zll_main_inputs_in[37:32], zll_main_inputs_in[31:15], zll_main_inputs_in[14:0]};
  assign zll_main_inputs6_in = {zll_main_inputs2_in[53:46], zll_main_inputs2_in[45:38], zll_main_inputs2_in[37:32], zll_main_inputs2_in[31:15], zll_main_inputs2_in[14:0]};
  assign zll_main_inputs3_in = {zll_main_inputs6_in[45:38], zll_main_inputs6_in[37:32], zll_main_inputs6_in[31:15], zll_main_inputs6_in[14:0]};
  assign zll_main_inputs1_in = {zll_main_inputs3_in[37:32], zll_main_inputs3_in[31:15], zll_main_inputs3_in[14:0]};
  assign zll_main_inputs4_in = {zll_main_inputs1_in[31:15], zll_main_inputs1_in[14:0]};
  assign res = {zll_main_inputs4_in[31:15], zll_main_getins_in[69:0]};
endmodule

module ZLL_Main_loop138 (input logic [142:0] arg0,
  output logic [142:0] res);
  logic [142:0] zll_main_loop251_in;
  logic [69:0] main_loop_in;
  logic [69:0] main_getinstr_in;
  logic [69:0] main_getins_in;
  logic [86:0] main_getins_out;
  logic [86:0] zll_main_getinstr1_in;
  logic [86:0] zll_main_getinstr2_in;
  logic [16:0] main_instrin_in;
  logic [16:0] zll_main_instrin_in;
  logic [78:0] zll_main_loop35_in;
  logic [78:0] zll_main_loop258_in;
  logic [142:0] zll_main_loop119_in;
  logic [142:0] zll_main_loop253_in;
  logic [78:0] zll_main_loop88_in;
  logic [139:0] zll_main_loop82_in;
  logic [139:0] zll_main_loop190_in;
  logic [151:0] zll_main_loop128_in;
  logic [151:0] zll_main_loop153_in;
  logic [148:0] zll_main_loop174_in;
  logic [78:0] zll_main_loop48_in;
  logic [75:0] zll_main_loop234_in;
  logic [75:0] zll_main_loop225_in;
  logic [69:0] zll_main_getreg13_in;
  logic [77:0] zll_main_getreg13_out;
  logic [83:0] zll_main_loop155_in;
  logic [83:0] zll_main_loop134_in;
  logic [15:0] binop_in;
  logic [15:0] binop_inR1;
  logic [76:0] zll_main_loop83_in;
  logic [75:0] zll_main_loop8_in;
  logic [75:0] main_putpc1_in;
  logic [69:0] main_putpc1_out;
  logic [70:0] zll_main_loop224_in;
  logic [69:0] main_incrpc_in;
  logic [69:0] main_incrpc_out;
  logic [69:0] zll_main_loop259_in;
  logic [142:0] zll_main_loop259_out;
  logic [142:0] zll_main_loop95_in;
  logic [142:0] zll_main_loop186_in;
  logic [69:0] zll_main_loop69_in;
  logic [69:0] main_getpc_in;
  logic [75:0] main_getpc_out;
  logic [75:0] zll_main_loop247_in;
  logic [69:0] zll_main_loop247_out;
  logic [69:0] zll_main_loop259_inR1;
  logic [142:0] zll_main_loop259_outR1;
  logic [142:0] zll_main_loop160_in;
  logic [142:0] zll_main_loop89_in;
  logic [69:0] zll_main_loop129_in;
  logic [69:0] main_getout_in;
  logic [84:0] main_getout_out;
  logic [84:0] zll_main_loop260_in;
  logic [142:0] zll_main_loop260_out;
  logic [142:0] zll_main_loop203_in;
  logic [142:0] zll_main_loop86_in;
  logic [84:0] zll_main_loop5_in;
  logic [78:0] zll_main_loop235_in;
  logic [75:0] zll_main_loop176_in;
  logic [75:0] zll_main_loop204_in;
  logic [71:0] main_getreg1_in;
  logic [77:0] main_getreg1_out;
  logic [81:0] zll_main_loop117_in;
  logic [81:0] zll_main_loop68_in;
  logic [81:0] zll_main_loop177_in;
  logic [71:0] main_getreg1_inR1;
  logic [77:0] main_getreg1_outR1;
  logic [87:0] zll_main_loop187_in;
  logic [87:0] zll_main_loop141_in;
  logic [15:0] binop_inR2;
  logic [7:0] unop_in;
  logic [79:0] main_putreg_in;
  logic [79:0] zll_main_putreg30_in;
  logic [77:0] zll_main_putreg43_in;
  logic [77:0] zll_main_putreg17_in;
  logic [147:0] zll_main_putreg8_in;
  logic [147:0] zll_main_putreg21_in;
  logic [77:0] zll_main_putreg31_in;
  logic [77:0] zll_main_putreg15_in;
  logic [79:0] zll_main_putreg28_in;
  logic [77:0] zll_main_putreg16_in;
  logic [77:0] zll_main_putreg22_in;
  logic [147:0] zll_main_putreg42_in;
  logic [147:0] zll_main_putreg2_in;
  logic [77:0] zll_main_putreg40_in;
  logic [79:0] zll_main_putreg20_in;
  logic [77:0] zll_main_putreg33_in;
  logic [77:0] zll_main_putreg9_in;
  logic [147:0] zll_main_putreg13_in;
  logic [147:0] zll_main_putreg7_in;
  logic [77:0] zll_main_putreg47_in;
  logic [79:0] zll_main_putreg5_in;
  logic [77:0] zll_main_putreg41_in;
  logic [77:0] main_putreg1_in;
  logic [69:0] main_putreg1_out;
  logic [69:0] main_incrpc_inR1;
  logic [69:0] main_incrpc_outR1;
  logic [69:0] zll_main_loop259_inR2;
  logic [142:0] zll_main_loop259_outR2;
  logic [142:0] zll_main_loop226_in;
  logic [142:0] zll_main_loop198_in;
  logic [69:0] zll_main_loop94_in;
  logic [69:0] main_getpc_inR1;
  logic [75:0] main_getpc_outR1;
  logic [75:0] zll_main_loop247_inR1;
  logic [69:0] zll_main_loop247_outR1;
  logic [69:0] zll_main_loop259_inR3;
  logic [142:0] zll_main_loop259_outR3;
  logic [142:0] zll_main_loop92_in;
  logic [142:0] zll_main_loop219_in;
  logic [69:0] zll_main_loop106_in;
  logic [69:0] main_getout_inR1;
  logic [84:0] main_getout_outR1;
  logic [84:0] zll_main_loop260_inR1;
  logic [142:0] zll_main_loop260_outR1;
  logic [142:0] zll_main_loop50_in;
  logic [142:0] zll_main_loop32_in;
  logic [84:0] zll_main_loop63_in;
  logic [78:0] zll_main_loop75_in;
  logic [75:0] zll_main_loop229_in;
  logic [75:0] zll_main_loop4_in;
  logic [69:0] zll_main_getreg13_inR1;
  logic [77:0] zll_main_getreg13_outR1;
  logic [83:0] zll_main_loop12_in;
  logic [83:0] zll_main_loop178_in;
  logic [75:0] main_putaddrout_in;
  logic [69:0] main_putaddrout_out;
  logic [77:0] zll_main_loop218_in;
  logic [77:0] main_putdataout1_in;
  logic [69:0] main_getout_inR2;
  logic [84:0] main_getout_outR2;
  logic [92:0] zll_main_putdataout2_in;
  logic [92:0] zll_main_putdataout8_in;
  logic [22:0] zll_main_putdataout_in;
  logic [22:0] zll_main_putdataout5_in;
  logic [22:0] zll_main_putdataout10_in;
  logic [84:0] main_putout_in;
  logic [69:0] main_putout_out;
  logic [69:0] main_putweout_in;
  logic [69:0] main_getout_inR3;
  logic [84:0] main_getout_outR3;
  logic [84:0] zll_main_putweout5_in;
  logic [84:0] zll_main_putweout2_in;
  logic [14:0] zll_main_putweout_in;
  logic [84:0] main_putout_inR1;
  logic [69:0] main_putout_outR1;
  logic [69:0] zll_main_loop259_inR4;
  logic [142:0] zll_main_loop259_outR4;
  logic [142:0] zll_main_loop74_in;
  logic [142:0] zll_main_loop216_in;
  logic [69:0] zll_main_loop154_in;
  logic [69:0] main_getout_inR4;
  logic [84:0] main_getout_outR4;
  logic [84:0] zll_main_loop260_inR2;
  logic [142:0] zll_main_loop260_outR2;
  logic [142:0] zll_main_loop209_in;
  logic [142:0] zll_main_loop236_in;
  logic [84:0] zll_main_loop81_in;
  logic [78:0] zll_main_loop256_in;
  logic [75:0] zll_main_loop64_in;
  logic [75:0] zll_main_loop77_in;
  logic [75:0] main_putaddrout_inR1;
  logic [69:0] main_putaddrout_outR1;
  logic [69:0] main_putweout1_in;
  logic [69:0] main_putweout1_out;
  logic [69:0] zll_main_loop259_inR5;
  logic [142:0] zll_main_loop259_outR5;
  logic [142:0] zll_main_loop113_in;
  logic [142:0] zll_main_loop205_in;
  logic [69:0] zll_main_loop118_in;
  logic [69:0] main_getout_inR5;
  logic [84:0] main_getout_outR5;
  logic [84:0] zll_main_loop260_inR3;
  logic [142:0] zll_main_loop260_outR3;
  logic [142:0] zll_main_loop151_in;
  logic [142:0] zll_main_loop212_in;
  logic [84:0] zll_main_loop150_in;
  logic [78:0] zll_main_loop242_in;
  logic [69:0] zll_main_loop175_in;
  logic [69:0] main_incrpc_inR2;
  logic [69:0] main_incrpc_outR2;
  logic [69:0] zll_main_loop259_inR6;
  logic [142:0] zll_main_loop259_outR6;
  logic [142:0] zll_main_loop170_in;
  logic [142:0] zll_main_loop15_in;
  logic [69:0] zll_main_loop228_in;
  logic [69:0] main_getpc_inR2;
  logic [75:0] main_getpc_outR2;
  logic [75:0] zll_main_loop247_inR2;
  logic [69:0] zll_main_loop247_outR2;
  logic [69:0] zll_main_loop259_inR7;
  logic [142:0] zll_main_loop259_outR7;
  logic [142:0] zll_main_loop45_in;
  logic [142:0] zll_main_loop241_in;
  logic [69:0] zll_main_loop139_in;
  logic [69:0] main_getout_inR6;
  logic [84:0] main_getout_outR6;
  logic [84:0] zll_main_loop260_inR4;
  logic [142:0] zll_main_loop260_outR4;
  logic [142:0] zll_main_loop91_in;
  logic [142:0] zll_main_loop98_in;
  logic [84:0] zll_main_loop231_in;
  assign zll_main_loop251_in = arg0;
  assign main_loop_in = zll_main_loop251_in[69:0];
  assign main_getinstr_in = main_loop_in[69:0];
  assign main_getins_in = main_getinstr_in[69:0];
  Main_getIns  inst (main_getins_in[69:0], main_getins_out);
  assign zll_main_getinstr1_in = main_getins_out;
  assign zll_main_getinstr2_in = zll_main_getinstr1_in[86:0];
  assign main_instrin_in = zll_main_getinstr2_in[86:70];
  assign zll_main_instrin_in = main_instrin_in[16:0];
  assign zll_main_loop35_in = {zll_main_instrin_in[16:8], zll_main_getinstr2_in[69:0]};
  assign zll_main_loop258_in = zll_main_loop35_in[78:0];
  assign zll_main_loop119_in = {{3'h1, {6'h3d{1'h0}}}, zll_main_loop258_in[78:70], zll_main_loop258_in[69:0]};
  assign zll_main_loop253_in = zll_main_loop119_in[142:0];
  assign zll_main_loop88_in = {zll_main_loop253_in[78:70], zll_main_loop253_in[69:0]};
  assign zll_main_loop82_in = {zll_main_loop88_in[69:0], zll_main_loop88_in[69:0]};
  assign zll_main_loop190_in = zll_main_loop82_in[139:0];
  assign zll_main_loop128_in = {zll_main_loop88_in[78:70], {3'h3, zll_main_loop190_in[139:70], zll_main_loop190_in[69:0]}};
  assign zll_main_loop153_in = {zll_main_loop128_in[151:143], zll_main_loop128_in[142:0]};
  assign zll_main_loop174_in = {zll_main_loop153_in[151:143], zll_main_loop153_in[139:70], zll_main_loop153_in[69:0]};
  assign zll_main_loop48_in = {zll_main_loop174_in[69:0], zll_main_loop174_in[148:140]};
  assign zll_main_loop234_in = {zll_main_loop48_in[78:9], zll_main_loop48_in[5:0]};
  assign zll_main_loop225_in = {zll_main_loop234_in[5:0], zll_main_loop234_in[75:6]};
  assign zll_main_getreg13_in = zll_main_loop225_in[69:0];
  ZLL_Main_getReg13  instR1 (zll_main_getreg13_in[69:0], zll_main_getreg13_out);
  assign zll_main_loop155_in = {zll_main_loop225_in[75:70], zll_main_getreg13_out};
  assign zll_main_loop134_in = {zll_main_loop155_in[83:78], zll_main_loop155_in[77:0]};
  assign binop_in = {zll_main_loop134_in[77:70], 8'h00};
  assign binop_inR1 = {zll_main_loop134_in[77:70], 8'h00};
  assign zll_main_loop83_in = {zll_main_loop134_in[69:0], zll_main_loop134_in[83:78], binop_inR1[15:8] == binop_inR1[7:0]};
  assign zll_main_loop8_in = {zll_main_loop83_in[76:7], zll_main_loop83_in[6:1]};
  assign main_putpc1_in = {zll_main_loop8_in[5:0], zll_main_loop8_in[75:6]};
  Main_putPC1  instR2 (main_putpc1_in[75:70], main_putpc1_in[69:0], main_putpc1_out);
  assign zll_main_loop224_in = {zll_main_loop134_in[69:0], binop_in[15:8] == binop_in[7:0]};
  assign main_incrpc_in = zll_main_loop224_in[70:1];
  Main_incrPC  instR3 (main_incrpc_in[69:0], main_incrpc_out);
  assign zll_main_loop259_in = (zll_main_loop224_in[0] == 1'h1) ? main_incrpc_out : main_putpc1_out;
  ZLL_Main_loop259  instR4 (zll_main_loop259_in[69:0], zll_main_loop259_out);
  assign zll_main_loop95_in = zll_main_loop259_out;
  assign zll_main_loop186_in = zll_main_loop95_in[142:0];
  assign zll_main_loop69_in = zll_main_loop186_in[69:0];
  assign main_getpc_in = zll_main_loop69_in[69:0];
  Main_getPC  instR5 (main_getpc_in[69:0], main_getpc_out);
  assign zll_main_loop247_in = main_getpc_out;
  ZLL_Main_loop247  instR6 (zll_main_loop247_in[75:0], zll_main_loop247_out);
  assign zll_main_loop259_inR1 = zll_main_loop247_out;
  ZLL_Main_loop259  instR7 (zll_main_loop259_inR1[69:0], zll_main_loop259_outR1);
  assign zll_main_loop160_in = zll_main_loop259_outR1;
  assign zll_main_loop89_in = zll_main_loop160_in[142:0];
  assign zll_main_loop129_in = zll_main_loop89_in[69:0];
  assign main_getout_in = zll_main_loop129_in[69:0];
  Main_getOut  instR8 (main_getout_in[69:0], main_getout_out);
  assign zll_main_loop260_in = main_getout_out;
  ZLL_Main_loop260  instR9 (zll_main_loop260_in[84:0], zll_main_loop260_out);
  assign zll_main_loop203_in = zll_main_loop260_out;
  assign zll_main_loop86_in = zll_main_loop203_in[142:0];
  assign zll_main_loop5_in = {zll_main_loop86_in[84:70], zll_main_loop86_in[69:0]};
  assign zll_main_loop235_in = {zll_main_loop174_in[69:0], zll_main_loop174_in[148:140]};
  assign zll_main_loop176_in = {zll_main_loop235_in[78:9], zll_main_loop235_in[5:4], zll_main_loop235_in[3:2], zll_main_loop235_in[1:0]};
  assign zll_main_loop204_in = {zll_main_loop176_in[5:4], zll_main_loop176_in[3:2], zll_main_loop176_in[1:0], zll_main_loop176_in[75:6]};
  assign main_getreg1_in = {zll_main_loop204_in[73:72], zll_main_loop204_in[69:0]};
  Main_getReg1  instR10 (main_getreg1_in[71:70], main_getreg1_in[69:0], main_getreg1_out);
  assign zll_main_loop117_in = {zll_main_loop204_in[75:74], zll_main_loop204_in[71:70], main_getreg1_out};
  assign zll_main_loop68_in = {zll_main_loop117_in[81:80], zll_main_loop117_in[79:78], zll_main_loop117_in[77:0]};
  assign zll_main_loop177_in = {zll_main_loop68_in[79:78], zll_main_loop68_in[81:80], zll_main_loop68_in[77:70], zll_main_loop68_in[69:0]};
  assign main_getreg1_inR1 = {zll_main_loop177_in[81:80], zll_main_loop177_in[69:0]};
  Main_getReg1  instR11 (main_getreg1_inR1[71:70], main_getreg1_inR1[69:0], main_getreg1_outR1);
  assign zll_main_loop187_in = {zll_main_loop177_in[79:78], zll_main_loop177_in[77:70], main_getreg1_outR1};
  assign zll_main_loop141_in = {zll_main_loop187_in[87:86], zll_main_loop187_in[85:78], zll_main_loop187_in[77:0]};
  assign binop_inR2 = {zll_main_loop141_in[85:78], zll_main_loop141_in[77:70]};
  assign unop_in = binop_inR2[15:8] & binop_inR2[7:0];
  assign main_putreg_in = {zll_main_loop141_in[87:86], ~unop_in[7:0], zll_main_loop141_in[69:0]};
  assign zll_main_putreg30_in = {main_putreg_in[69:0], main_putreg_in[79:78], main_putreg_in[77:70]};
  assign zll_main_putreg43_in = {zll_main_putreg30_in[79:10], zll_main_putreg30_in[7:0]};
  assign zll_main_putreg17_in = {zll_main_putreg43_in[7:0], zll_main_putreg43_in[77:8]};
  assign zll_main_putreg8_in = {zll_main_putreg17_in[77:70], zll_main_putreg17_in[69:0], zll_main_putreg17_in[69:0]};
  assign zll_main_putreg21_in = {zll_main_putreg8_in[147:140], zll_main_putreg8_in[139:0]};
  assign zll_main_putreg31_in = {zll_main_putreg21_in[147:140], zll_main_putreg21_in[139:70]};
  assign zll_main_putreg15_in = {zll_main_putreg31_in[61:54], zll_main_putreg31_in[77:70], zll_main_putreg31_in[69:62], zll_main_putreg31_in[53:46], zll_main_putreg31_in[45:38], zll_main_putreg31_in[37:32], zll_main_putreg31_in[31:15], zll_main_putreg31_in[14:0]};
  assign zll_main_putreg28_in = {main_putreg_in[69:0], main_putreg_in[79:78], main_putreg_in[77:70]};
  assign zll_main_putreg16_in = {zll_main_putreg28_in[79:10], zll_main_putreg28_in[7:0]};
  assign zll_main_putreg22_in = {zll_main_putreg16_in[7:0], zll_main_putreg16_in[77:8]};
  assign zll_main_putreg42_in = {zll_main_putreg22_in[77:70], zll_main_putreg22_in[69:0], zll_main_putreg22_in[69:0]};
  assign zll_main_putreg2_in = {zll_main_putreg42_in[147:140], zll_main_putreg42_in[139:0]};
  assign zll_main_putreg40_in = {zll_main_putreg2_in[147:140], zll_main_putreg2_in[139:70]};
  assign zll_main_putreg20_in = {main_putreg_in[69:0], main_putreg_in[79:78], main_putreg_in[77:70]};
  assign zll_main_putreg33_in = {zll_main_putreg20_in[79:10], zll_main_putreg20_in[7:0]};
  assign zll_main_putreg9_in = {zll_main_putreg33_in[7:0], zll_main_putreg33_in[77:8]};
  assign zll_main_putreg13_in = {zll_main_putreg9_in[77:70], zll_main_putreg9_in[69:0], zll_main_putreg9_in[69:0]};
  assign zll_main_putreg7_in = {zll_main_putreg13_in[147:140], zll_main_putreg13_in[139:0]};
  assign zll_main_putreg47_in = {zll_main_putreg7_in[147:140], zll_main_putreg7_in[139:70]};
  assign zll_main_putreg5_in = {main_putreg_in[69:0], main_putreg_in[79:78], main_putreg_in[77:70]};
  assign zll_main_putreg41_in = {zll_main_putreg5_in[79:10], zll_main_putreg5_in[7:0]};
  assign main_putreg1_in = {zll_main_putreg41_in[7:0], zll_main_putreg41_in[77:8]};
  Main_putReg1  instR12 (main_putreg1_in[77:70], main_putreg1_in[69:0], main_putreg1_out);
  assign main_incrpc_inR1 = (zll_main_putreg5_in[9:8] == 2'h0) ? main_putreg1_out : ((zll_main_putreg20_in[9:8] == 2'h1) ? {zll_main_putreg47_in[69:62], zll_main_putreg47_in[77:70], zll_main_putreg47_in[53:46], zll_main_putreg47_in[45:38], zll_main_putreg47_in[37:32], zll_main_putreg47_in[31:15], zll_main_putreg47_in[14:0]} : ((zll_main_putreg28_in[9:8] == 2'h2) ? {zll_main_putreg40_in[69:62], zll_main_putreg40_in[61:54], zll_main_putreg40_in[77:70], zll_main_putreg40_in[45:38], zll_main_putreg40_in[37:32], zll_main_putreg40_in[31:15], zll_main_putreg40_in[14:0]} : {zll_main_putreg15_in[61:54], zll_main_putreg15_in[77:70], zll_main_putreg15_in[53:46], zll_main_putreg15_in[69:62], zll_main_putreg15_in[37:32], zll_main_putreg15_in[31:15], zll_main_putreg15_in[14:0]}));
  Main_incrPC  instR13 (main_incrpc_inR1[69:0], main_incrpc_outR1);
  assign zll_main_loop259_inR2 = main_incrpc_outR1;
  ZLL_Main_loop259  instR14 (zll_main_loop259_inR2[69:0], zll_main_loop259_outR2);
  assign zll_main_loop226_in = zll_main_loop259_outR2;
  assign zll_main_loop198_in = zll_main_loop226_in[142:0];
  assign zll_main_loop94_in = zll_main_loop198_in[69:0];
  assign main_getpc_inR1 = zll_main_loop94_in[69:0];
  Main_getPC  instR15 (main_getpc_inR1[69:0], main_getpc_outR1);
  assign zll_main_loop247_inR1 = main_getpc_outR1;
  ZLL_Main_loop247  instR16 (zll_main_loop247_inR1[75:0], zll_main_loop247_outR1);
  assign zll_main_loop259_inR3 = zll_main_loop247_outR1;
  ZLL_Main_loop259  instR17 (zll_main_loop259_inR3[69:0], zll_main_loop259_outR3);
  assign zll_main_loop92_in = zll_main_loop259_outR3;
  assign zll_main_loop219_in = zll_main_loop92_in[142:0];
  assign zll_main_loop106_in = zll_main_loop219_in[69:0];
  assign main_getout_inR1 = zll_main_loop106_in[69:0];
  Main_getOut  instR18 (main_getout_inR1[69:0], main_getout_outR1);
  assign zll_main_loop260_inR1 = main_getout_outR1;
  ZLL_Main_loop260  instR19 (zll_main_loop260_inR1[84:0], zll_main_loop260_outR1);
  assign zll_main_loop50_in = zll_main_loop260_outR1;
  assign zll_main_loop32_in = zll_main_loop50_in[142:0];
  assign zll_main_loop63_in = {zll_main_loop32_in[84:70], zll_main_loop32_in[69:0]};
  assign zll_main_loop75_in = {zll_main_loop174_in[69:0], zll_main_loop174_in[148:140]};
  assign zll_main_loop229_in = {zll_main_loop75_in[78:9], zll_main_loop75_in[5:0]};
  assign zll_main_loop4_in = {zll_main_loop229_in[5:0], zll_main_loop229_in[75:6]};
  assign zll_main_getreg13_inR1 = zll_main_loop4_in[69:0];
  ZLL_Main_getReg13  instR20 (zll_main_getreg13_inR1[69:0], zll_main_getreg13_outR1);
  assign zll_main_loop12_in = {zll_main_loop4_in[75:70], zll_main_getreg13_outR1};
  assign zll_main_loop178_in = {zll_main_loop12_in[83:78], zll_main_loop12_in[77:0]};
  assign main_putaddrout_in = {zll_main_loop178_in[83:78], zll_main_loop178_in[69:0]};
  Main_putAddrOut  instR21 (main_putaddrout_in[75:70], main_putaddrout_in[69:0], main_putaddrout_out);
  assign zll_main_loop218_in = {zll_main_loop178_in[77:70], main_putaddrout_out};
  assign main_putdataout1_in = {zll_main_loop218_in[77:70], zll_main_loop218_in[69:0]};
  assign main_getout_inR2 = main_putdataout1_in[69:0];
  Main_getOut  instR22 (main_getout_inR2[69:0], main_getout_outR2);
  assign zll_main_putdataout2_in = {main_putdataout1_in[77:70], main_getout_outR2};
  assign zll_main_putdataout8_in = {zll_main_putdataout2_in[92:85], zll_main_putdataout2_in[84:0]};
  assign zll_main_putdataout_in = {zll_main_putdataout8_in[92:85], zll_main_putdataout8_in[84:70]};
  assign zll_main_putdataout5_in = {zll_main_putdataout_in[14], zll_main_putdataout_in[22:15], zll_main_putdataout_in[13:8], zll_main_putdataout_in[7:0]};
  assign zll_main_putdataout10_in = {zll_main_putdataout5_in[13:8], zll_main_putdataout5_in[22], zll_main_putdataout5_in[21:14], zll_main_putdataout5_in[7:0]};
  assign main_putout_in = {{zll_main_putdataout10_in[16], zll_main_putdataout10_in[22:17], zll_main_putdataout10_in[15:8]}, zll_main_putdataout8_in[69:0]};
  Main_putOut  instR23 (main_putout_in[84:70], main_putout_in[69:0], main_putout_out);
  assign main_putweout_in = main_putout_out;
  assign main_getout_inR3 = main_putweout_in[69:0];
  Main_getOut  instR24 (main_getout_inR3[69:0], main_getout_outR3);
  assign zll_main_putweout5_in = main_getout_outR3;
  assign zll_main_putweout2_in = zll_main_putweout5_in[84:0];
  assign zll_main_putweout_in = zll_main_putweout2_in[84:70];
  assign main_putout_inR1 = {{1'h1, zll_main_putweout_in[13:8], zll_main_putweout_in[7:0]}, zll_main_putweout2_in[69:0]};
  Main_putOut  instR25 (main_putout_inR1[84:70], main_putout_inR1[69:0], main_putout_outR1);
  assign zll_main_loop259_inR4 = main_putout_outR1;
  ZLL_Main_loop259  instR26 (zll_main_loop259_inR4[69:0], zll_main_loop259_outR4);
  assign zll_main_loop74_in = zll_main_loop259_outR4;
  assign zll_main_loop216_in = zll_main_loop74_in[142:0];
  assign zll_main_loop154_in = zll_main_loop216_in[69:0];
  assign main_getout_inR4 = zll_main_loop154_in[69:0];
  Main_getOut  instR27 (main_getout_inR4[69:0], main_getout_outR4);
  assign zll_main_loop260_inR2 = main_getout_outR4;
  ZLL_Main_loop260  instR28 (zll_main_loop260_inR2[84:0], zll_main_loop260_outR2);
  assign zll_main_loop209_in = zll_main_loop260_outR2;
  assign zll_main_loop236_in = zll_main_loop209_in[142:0];
  assign zll_main_loop81_in = {zll_main_loop236_in[84:70], zll_main_loop236_in[69:0]};
  assign zll_main_loop256_in = {zll_main_loop174_in[69:0], zll_main_loop174_in[148:140]};
  assign zll_main_loop64_in = {zll_main_loop256_in[78:9], zll_main_loop256_in[5:0]};
  assign zll_main_loop77_in = {zll_main_loop64_in[5:0], zll_main_loop64_in[75:6]};
  assign main_putaddrout_inR1 = {zll_main_loop77_in[75:70], zll_main_loop77_in[69:0]};
  Main_putAddrOut  instR29 (main_putaddrout_inR1[75:70], main_putaddrout_inR1[69:0], main_putaddrout_outR1);
  assign main_putweout1_in = main_putaddrout_outR1;
  Main_putWeOut1  instR30 (main_putweout1_in[69:0], main_putweout1_out);
  assign zll_main_loop259_inR5 = main_putweout1_out;
  ZLL_Main_loop259  instR31 (zll_main_loop259_inR5[69:0], zll_main_loop259_outR5);
  assign zll_main_loop113_in = zll_main_loop259_outR5;
  assign zll_main_loop205_in = zll_main_loop113_in[142:0];
  assign zll_main_loop118_in = zll_main_loop205_in[69:0];
  assign main_getout_inR5 = zll_main_loop118_in[69:0];
  Main_getOut  instR32 (main_getout_inR5[69:0], main_getout_outR5);
  assign zll_main_loop260_inR3 = main_getout_outR5;
  ZLL_Main_loop260  instR33 (zll_main_loop260_inR3[84:0], zll_main_loop260_outR3);
  assign zll_main_loop151_in = zll_main_loop260_outR3;
  assign zll_main_loop212_in = zll_main_loop151_in[142:0];
  assign zll_main_loop150_in = {zll_main_loop212_in[84:70], zll_main_loop212_in[69:0]};
  assign zll_main_loop242_in = {zll_main_loop174_in[69:0], zll_main_loop174_in[148:140]};
  assign zll_main_loop175_in = zll_main_loop242_in[78:9];
  assign main_incrpc_inR2 = zll_main_loop175_in[69:0];
  Main_incrPC  instR34 (main_incrpc_inR2[69:0], main_incrpc_outR2);
  assign zll_main_loop259_inR6 = main_incrpc_outR2;
  ZLL_Main_loop259  instR35 (zll_main_loop259_inR6[69:0], zll_main_loop259_outR6);
  assign zll_main_loop170_in = zll_main_loop259_outR6;
  assign zll_main_loop15_in = zll_main_loop170_in[142:0];
  assign zll_main_loop228_in = zll_main_loop15_in[69:0];
  assign main_getpc_inR2 = zll_main_loop228_in[69:0];
  Main_getPC  instR36 (main_getpc_inR2[69:0], main_getpc_outR2);
  assign zll_main_loop247_inR2 = main_getpc_outR2;
  ZLL_Main_loop247  instR37 (zll_main_loop247_inR2[75:0], zll_main_loop247_outR2);
  assign zll_main_loop259_inR7 = zll_main_loop247_outR2;
  ZLL_Main_loop259  instR38 (zll_main_loop259_inR7[69:0], zll_main_loop259_outR7);
  assign zll_main_loop45_in = zll_main_loop259_outR7;
  assign zll_main_loop241_in = zll_main_loop45_in[142:0];
  assign zll_main_loop139_in = zll_main_loop241_in[69:0];
  assign main_getout_inR6 = zll_main_loop139_in[69:0];
  Main_getOut  instR39 (main_getout_inR6[69:0], main_getout_outR6);
  assign zll_main_loop260_inR4 = main_getout_outR6;
  ZLL_Main_loop260  instR40 (zll_main_loop260_inR4[84:0], zll_main_loop260_outR4);
  assign zll_main_loop91_in = zll_main_loop260_outR4;
  assign zll_main_loop98_in = zll_main_loop91_in[142:0];
  assign zll_main_loop231_in = {zll_main_loop98_in[84:70], zll_main_loop98_in[69:0]};
  assign res = (zll_main_loop242_in[8:6] == 3'h0) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop231_in[84:70], 4'h0, zll_main_loop231_in[69:0]} : ((zll_main_loop256_in[8:6] == 3'h1) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop150_in[84:70], 4'h2, zll_main_loop150_in[69:0]} : ((zll_main_loop75_in[8:6] == 3'h2) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop81_in[84:70], 4'h4, zll_main_loop81_in[69:0]} : ((zll_main_loop235_in[8:6] == 3'h3) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop63_in[84:70], 4'h5, zll_main_loop63_in[69:0]} : {{1'h1, {6'h35{1'h0}}}, zll_main_loop5_in[84:70], 4'h6, zll_main_loop5_in[69:0]})));
endmodule

module Main_getOut (input logic [69:0] arg0,
  output logic [84:0] res);
  logic [139:0] zll_main_getout_in;
  logic [139:0] zll_main_getout1_in;
  logic [69:0] main_outputs_in;
  logic [69:0] zll_main_outputs2_in;
  logic [61:0] zll_main_outputs1_in;
  logic [53:0] zll_main_outputs3_in;
  logic [45:0] zll_main_outputs6_in;
  logic [37:0] zll_main_outputs5_in;
  logic [31:0] zll_main_outputs_in;
  assign zll_main_getout_in = {arg0, arg0};
  assign zll_main_getout1_in = zll_main_getout_in[139:0];
  assign main_outputs_in = zll_main_getout1_in[139:70];
  assign zll_main_outputs2_in = main_outputs_in[69:0];
  assign zll_main_outputs1_in = {zll_main_outputs2_in[61:54], zll_main_outputs2_in[53:46], zll_main_outputs2_in[45:38], zll_main_outputs2_in[37:32], zll_main_outputs2_in[31:15], zll_main_outputs2_in[14:0]};
  assign zll_main_outputs3_in = {zll_main_outputs1_in[53:46], zll_main_outputs1_in[45:38], zll_main_outputs1_in[37:32], zll_main_outputs1_in[31:15], zll_main_outputs1_in[14:0]};
  assign zll_main_outputs6_in = {zll_main_outputs3_in[45:38], zll_main_outputs3_in[37:32], zll_main_outputs3_in[31:15], zll_main_outputs3_in[14:0]};
  assign zll_main_outputs5_in = {zll_main_outputs6_in[37:32], zll_main_outputs6_in[31:15], zll_main_outputs6_in[14:0]};
  assign zll_main_outputs_in = {zll_main_outputs5_in[31:15], zll_main_outputs5_in[14:0]};
  assign res = {zll_main_outputs_in[14:0], zll_main_getout1_in[69:0]};
endmodule

module Main_putAddrOut (input logic [5:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [69:0] main_getout_in;
  logic [84:0] main_getout_out;
  logic [90:0] zll_main_putaddrout6_in;
  logic [90:0] zll_main_putaddrout_in;
  logic [20:0] zll_main_putaddrout4_in;
  logic [20:0] zll_main_putaddrout5_in;
  logic [84:0] main_putout_in;
  logic [69:0] main_putout_out;
  assign main_getout_in = arg1;
  Main_getOut  inst (main_getout_in[69:0], main_getout_out);
  assign zll_main_putaddrout6_in = {arg0, main_getout_out};
  assign zll_main_putaddrout_in = {zll_main_putaddrout6_in[90:85], zll_main_putaddrout6_in[84:0]};
  assign zll_main_putaddrout4_in = {zll_main_putaddrout_in[90:85], zll_main_putaddrout_in[84:70]};
  assign zll_main_putaddrout5_in = {zll_main_putaddrout4_in[14], zll_main_putaddrout4_in[20:15], zll_main_putaddrout4_in[13:8], zll_main_putaddrout4_in[7:0]};
  assign main_putout_in = {{zll_main_putaddrout5_in[20], zll_main_putaddrout5_in[19:14], zll_main_putaddrout5_in[7:0]}, zll_main_putaddrout_in[69:0]};
  Main_putOut  instR1 (main_putout_in[84:70], main_putout_in[69:0], main_putout_out);
  assign res = main_putout_out;
endmodule

module Main_incrPC (input logic [69:0] arg0,
  output logic [69:0] res);
  logic [69:0] main_getpc_in;
  logic [75:0] main_getpc_out;
  logic [75:0] zll_main_incrpc1_in;
  logic [75:0] zll_main_incrpc_in;
  logic [11:0] binop_in;
  logic [75:0] main_putpc1_in;
  logic [69:0] main_putpc1_out;
  assign main_getpc_in = arg0;
  Main_getPC  inst (main_getpc_in[69:0], main_getpc_out);
  assign zll_main_incrpc1_in = main_getpc_out;
  assign zll_main_incrpc_in = zll_main_incrpc1_in[75:0];
  assign binop_in = {zll_main_incrpc_in[75:70], 6'h01};
  assign main_putpc1_in = {binop_in[11:6] + binop_in[5:0], zll_main_incrpc_in[69:0]};
  Main_putPC1  instR1 (main_putpc1_in[75:70], main_putpc1_in[69:0], main_putpc1_out);
  assign res = main_putpc1_out;
endmodule

module Main_getPC (input logic [69:0] arg0,
  output logic [75:0] res);
  logic [139:0] zll_main_getpc_in;
  logic [139:0] zll_main_getpc1_in;
  logic [69:0] main_pc_in;
  logic [69:0] zll_main_pc5_in;
  logic [61:0] zll_main_pc4_in;
  logic [53:0] zll_main_pc_in;
  logic [45:0] zll_main_pc6_in;
  logic [37:0] zll_main_pc3_in;
  logic [20:0] zll_main_pc2_in;
  assign zll_main_getpc_in = {arg0, arg0};
  assign zll_main_getpc1_in = zll_main_getpc_in[139:0];
  assign main_pc_in = zll_main_getpc1_in[139:70];
  assign zll_main_pc5_in = main_pc_in[69:0];
  assign zll_main_pc4_in = {zll_main_pc5_in[61:54], zll_main_pc5_in[53:46], zll_main_pc5_in[45:38], zll_main_pc5_in[37:32], zll_main_pc5_in[31:15], zll_main_pc5_in[14:0]};
  assign zll_main_pc_in = {zll_main_pc4_in[53:46], zll_main_pc4_in[45:38], zll_main_pc4_in[37:32], zll_main_pc4_in[31:15], zll_main_pc4_in[14:0]};
  assign zll_main_pc6_in = {zll_main_pc_in[45:38], zll_main_pc_in[37:32], zll_main_pc_in[31:15], zll_main_pc_in[14:0]};
  assign zll_main_pc3_in = {zll_main_pc6_in[37:32], zll_main_pc6_in[31:15], zll_main_pc6_in[14:0]};
  assign zll_main_pc2_in = {zll_main_pc3_in[37:32], zll_main_pc3_in[14:0]};
  assign res = {zll_main_pc2_in[20:15], zll_main_getpc1_in[69:0]};
endmodule

module Main_putOut (input logic [14:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [154:0] zll_main_putout3_in;
  logic [154:0] zll_main_putout11_in;
  logic [84:0] zll_main_putout5_in;
  logic [84:0] zll_main_putout8_in;
  logic [84:0] zll_main_putout9_in;
  assign zll_main_putout3_in = {arg0, arg1, arg1};
  assign zll_main_putout11_in = {zll_main_putout3_in[154:140], zll_main_putout3_in[139:0]};
  assign zll_main_putout5_in = {zll_main_putout11_in[154:140], zll_main_putout11_in[139:70]};
  assign zll_main_putout8_in = {zll_main_putout5_in[53:46], zll_main_putout5_in[84:70], zll_main_putout5_in[69:62], zll_main_putout5_in[61:54], zll_main_putout5_in[45:38], zll_main_putout5_in[37:32], zll_main_putout5_in[31:15], zll_main_putout5_in[14:0]};
  assign zll_main_putout9_in = {zll_main_putout8_in[84:77], zll_main_putout8_in[31:15], zll_main_putout8_in[76:62], zll_main_putout8_in[61:54], zll_main_putout8_in[53:46], zll_main_putout8_in[45:38], zll_main_putout8_in[37:32], zll_main_putout8_in[14:0]};
  assign res = {zll_main_putout9_in[44:37], zll_main_putout9_in[36:29], zll_main_putout9_in[84:77], zll_main_putout9_in[28:21], zll_main_putout9_in[20:15], zll_main_putout9_in[76:60], zll_main_putout9_in[59:45]};
endmodule