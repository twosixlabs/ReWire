module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [99:0] __in0,
  output logic [99:0] __out0,
  output logic [99:0] __out1,
  output logic [99:0] __out2,
  output logic [99:0] __out3);
  logic [99:0] gMainzidev;
  logic [106:0] gzdLLziMainzidev2;
  logic [0:0] callRes;
  logic [106:0] gzdLLziMainzidev2R1;
  logic [0:0] callResR1;
  logic [106:0] gzdLLziMainzidev2R2;
  logic [0:0] callResR2;
  logic [106:0] gzdLLziMainzidev2R3;
  logic [0:0] callResR3;
  logic [106:0] gzdLLziMainzidev2R4;
  logic [0:0] callResR4;
  logic [106:0] gzdLLziMainzidev2R5;
  logic [0:0] callResR5;
  logic [106:0] gzdLLziMainzidev2R6;
  logic [0:0] callResR6;
  logic [106:0] gzdLLziMainzidev2R7;
  logic [0:0] callResR7;
  logic [106:0] gzdLLziMainzidev2R8;
  logic [0:0] callResR8;
  logic [106:0] gzdLLziMainzidev2R9;
  logic [0:0] callResR9;
  logic [106:0] gzdLLziMainzidev2R10;
  logic [0:0] callResR10;
  logic [106:0] gzdLLziMainzidev2R11;
  logic [0:0] callResR11;
  logic [106:0] gzdLLziMainzidev2R12;
  logic [0:0] callResR12;
  logic [106:0] gzdLLziMainzidev2R13;
  logic [0:0] callResR13;
  logic [106:0] gzdLLziMainzidev2R14;
  logic [0:0] callResR14;
  logic [106:0] gzdLLziMainzidev2R15;
  logic [0:0] callResR15;
  logic [106:0] gzdLLziMainzidev2R16;
  logic [0:0] callResR16;
  logic [106:0] gzdLLziMainzidev2R17;
  logic [0:0] callResR17;
  logic [106:0] gzdLLziMainzidev2R18;
  logic [0:0] callResR18;
  logic [106:0] gzdLLziMainzidev2R19;
  logic [0:0] callResR19;
  logic [106:0] gzdLLziMainzidev2R20;
  logic [0:0] callResR20;
  logic [106:0] gzdLLziMainzidev2R21;
  logic [0:0] callResR21;
  logic [106:0] gzdLLziMainzidev2R22;
  logic [0:0] callResR22;
  logic [106:0] gzdLLziMainzidev2R23;
  logic [0:0] callResR23;
  logic [106:0] gzdLLziMainzidev2R24;
  logic [0:0] callResR24;
  logic [106:0] gzdLLziMainzidev2R25;
  logic [0:0] callResR25;
  logic [106:0] gzdLLziMainzidev2R26;
  logic [0:0] callResR26;
  logic [106:0] gzdLLziMainzidev2R27;
  logic [0:0] callResR27;
  logic [106:0] gzdLLziMainzidev2R28;
  logic [0:0] callResR28;
  logic [106:0] gzdLLziMainzidev2R29;
  logic [0:0] callResR29;
  logic [106:0] gzdLLziMainzidev2R30;
  logic [0:0] callResR30;
  logic [106:0] gzdLLziMainzidev2R31;
  logic [0:0] callResR31;
  logic [106:0] gzdLLziMainzidev2R32;
  logic [0:0] callResR32;
  logic [106:0] gzdLLziMainzidev2R33;
  logic [0:0] callResR33;
  logic [106:0] gzdLLziMainzidev2R34;
  logic [0:0] callResR34;
  logic [106:0] gzdLLziMainzidev2R35;
  logic [0:0] callResR35;
  logic [106:0] gzdLLziMainzidev2R36;
  logic [0:0] callResR36;
  logic [106:0] gzdLLziMainzidev2R37;
  logic [0:0] callResR37;
  logic [106:0] gzdLLziMainzidev2R38;
  logic [0:0] callResR38;
  logic [106:0] gzdLLziMainzidev2R39;
  logic [0:0] callResR39;
  logic [106:0] gzdLLziMainzidev2R40;
  logic [0:0] callResR40;
  logic [106:0] gzdLLziMainzidev2R41;
  logic [0:0] callResR41;
  logic [106:0] gzdLLziMainzidev2R42;
  logic [0:0] callResR42;
  logic [106:0] gzdLLziMainzidev2R43;
  logic [0:0] callResR43;
  logic [106:0] gzdLLziMainzidev2R44;
  logic [0:0] callResR44;
  logic [106:0] gzdLLziMainzidev2R45;
  logic [0:0] callResR45;
  logic [106:0] gzdLLziMainzidev2R46;
  logic [0:0] callResR46;
  logic [106:0] gzdLLziMainzidev2R47;
  logic [0:0] callResR47;
  logic [106:0] gzdLLziMainzidev2R48;
  logic [0:0] callResR48;
  logic [106:0] gzdLLziMainzidev2R49;
  logic [0:0] callResR49;
  logic [106:0] gzdLLziMainzidev2R50;
  logic [0:0] callResR50;
  logic [106:0] gzdLLziMainzidev2R51;
  logic [0:0] callResR51;
  logic [106:0] gzdLLziMainzidev2R52;
  logic [0:0] callResR52;
  logic [106:0] gzdLLziMainzidev2R53;
  logic [0:0] callResR53;
  logic [106:0] gzdLLziMainzidev2R54;
  logic [0:0] callResR54;
  logic [106:0] gzdLLziMainzidev2R55;
  logic [0:0] callResR55;
  logic [106:0] gzdLLziMainzidev2R56;
  logic [0:0] callResR56;
  logic [106:0] gzdLLziMainzidev2R57;
  logic [0:0] callResR57;
  logic [106:0] gzdLLziMainzidev2R58;
  logic [0:0] callResR58;
  logic [106:0] gzdLLziMainzidev2R59;
  logic [0:0] callResR59;
  logic [106:0] gzdLLziMainzidev2R60;
  logic [0:0] callResR60;
  logic [106:0] gzdLLziMainzidev2R61;
  logic [0:0] callResR61;
  logic [106:0] gzdLLziMainzidev2R62;
  logic [0:0] callResR62;
  logic [106:0] gzdLLziMainzidev2R63;
  logic [0:0] callResR63;
  logic [106:0] gzdLLziMainzidev2R64;
  logic [0:0] callResR64;
  logic [106:0] gzdLLziMainzidev2R65;
  logic [0:0] callResR65;
  logic [106:0] gzdLLziMainzidev2R66;
  logic [0:0] callResR66;
  logic [106:0] gzdLLziMainzidev2R67;
  logic [0:0] callResR67;
  logic [106:0] gzdLLziMainzidev2R68;
  logic [0:0] callResR68;
  logic [106:0] gzdLLziMainzidev2R69;
  logic [0:0] callResR69;
  logic [106:0] gzdLLziMainzidev2R70;
  logic [0:0] callResR70;
  logic [106:0] gzdLLziMainzidev2R71;
  logic [0:0] callResR71;
  logic [106:0] gzdLLziMainzidev2R72;
  logic [0:0] callResR72;
  logic [106:0] gzdLLziMainzidev2R73;
  logic [0:0] callResR73;
  logic [106:0] gzdLLziMainzidev2R74;
  logic [0:0] callResR74;
  logic [106:0] gzdLLziMainzidev2R75;
  logic [0:0] callResR75;
  logic [106:0] gzdLLziMainzidev2R76;
  logic [0:0] callResR76;
  logic [106:0] gzdLLziMainzidev2R77;
  logic [0:0] callResR77;
  logic [106:0] gzdLLziMainzidev2R78;
  logic [0:0] callResR78;
  logic [106:0] gzdLLziMainzidev2R79;
  logic [0:0] callResR79;
  logic [106:0] gzdLLziMainzidev2R80;
  logic [0:0] callResR80;
  logic [106:0] gzdLLziMainzidev2R81;
  logic [0:0] callResR81;
  logic [106:0] gzdLLziMainzidev2R82;
  logic [0:0] callResR82;
  logic [106:0] gzdLLziMainzidev2R83;
  logic [0:0] callResR83;
  logic [106:0] gzdLLziMainzidev2R84;
  logic [0:0] callResR84;
  logic [106:0] gzdLLziMainzidev2R85;
  logic [0:0] callResR85;
  logic [106:0] gzdLLziMainzidev2R86;
  logic [0:0] callResR86;
  logic [106:0] gzdLLziMainzidev2R87;
  logic [0:0] callResR87;
  logic [106:0] gzdLLziMainzidev2R88;
  logic [0:0] callResR88;
  logic [106:0] gzdLLziMainzidev2R89;
  logic [0:0] callResR89;
  logic [106:0] gzdLLziMainzidev2R90;
  logic [0:0] callResR90;
  logic [106:0] gzdLLziMainzidev2R91;
  logic [0:0] callResR91;
  logic [106:0] gzdLLziMainzidev2R92;
  logic [0:0] callResR92;
  logic [106:0] gzdLLziMainzidev2R93;
  logic [0:0] callResR93;
  logic [106:0] gzdLLziMainzidev2R94;
  logic [0:0] callResR94;
  logic [106:0] gzdLLziMainzidev2R95;
  logic [0:0] callResR95;
  logic [106:0] gzdLLziMainzidev2R96;
  logic [0:0] callResR96;
  logic [106:0] gzdLLziMainzidev2R97;
  logic [0:0] callResR97;
  logic [106:0] gzdLLziMainzidev2R98;
  logic [0:0] callResR98;
  logic [106:0] gzdLLziMainzidev2R99;
  logic [0:0] callResR99;
  logic [106:0] gzdLLziMainzidev5;
  logic [0:0] callResR100;
  logic [106:0] gzdLLziMainzidev5R1;
  logic [0:0] callResR101;
  logic [106:0] gzdLLziMainzidev5R2;
  logic [0:0] callResR102;
  logic [106:0] gzdLLziMainzidev5R3;
  logic [0:0] callResR103;
  logic [106:0] gzdLLziMainzidev5R4;
  logic [0:0] callResR104;
  logic [106:0] gzdLLziMainzidev5R5;
  logic [0:0] callResR105;
  logic [106:0] gzdLLziMainzidev5R6;
  logic [0:0] callResR106;
  logic [106:0] gzdLLziMainzidev5R7;
  logic [0:0] callResR107;
  logic [106:0] gzdLLziMainzidev5R8;
  logic [0:0] callResR108;
  logic [106:0] gzdLLziMainzidev5R9;
  logic [0:0] callResR109;
  logic [106:0] gzdLLziMainzidev5R10;
  logic [0:0] callResR110;
  logic [106:0] gzdLLziMainzidev5R11;
  logic [0:0] callResR111;
  logic [106:0] gzdLLziMainzidev5R12;
  logic [0:0] callResR112;
  logic [106:0] gzdLLziMainzidev5R13;
  logic [0:0] callResR113;
  logic [106:0] gzdLLziMainzidev5R14;
  logic [0:0] callResR114;
  logic [106:0] gzdLLziMainzidev5R15;
  logic [0:0] callResR115;
  logic [106:0] gzdLLziMainzidev5R16;
  logic [0:0] callResR116;
  logic [106:0] gzdLLziMainzidev5R17;
  logic [0:0] callResR117;
  logic [106:0] gzdLLziMainzidev5R18;
  logic [0:0] callResR118;
  logic [106:0] gzdLLziMainzidev5R19;
  logic [0:0] callResR119;
  logic [106:0] gzdLLziMainzidev5R20;
  logic [0:0] callResR120;
  logic [106:0] gzdLLziMainzidev5R21;
  logic [0:0] callResR121;
  logic [106:0] gzdLLziMainzidev5R22;
  logic [0:0] callResR122;
  logic [106:0] gzdLLziMainzidev5R23;
  logic [0:0] callResR123;
  logic [106:0] gzdLLziMainzidev5R24;
  logic [0:0] callResR124;
  logic [106:0] gzdLLziMainzidev5R25;
  logic [0:0] callResR125;
  logic [106:0] gzdLLziMainzidev5R26;
  logic [0:0] callResR126;
  logic [106:0] gzdLLziMainzidev5R27;
  logic [0:0] callResR127;
  logic [106:0] gzdLLziMainzidev5R28;
  logic [0:0] callResR128;
  logic [106:0] gzdLLziMainzidev5R29;
  logic [0:0] callResR129;
  logic [106:0] gzdLLziMainzidev5R30;
  logic [0:0] callResR130;
  logic [106:0] gzdLLziMainzidev5R31;
  logic [0:0] callResR131;
  logic [106:0] gzdLLziMainzidev5R32;
  logic [0:0] callResR132;
  logic [106:0] gzdLLziMainzidev5R33;
  logic [0:0] callResR133;
  logic [106:0] gzdLLziMainzidev5R34;
  logic [0:0] callResR134;
  logic [106:0] gzdLLziMainzidev5R35;
  logic [0:0] callResR135;
  logic [106:0] gzdLLziMainzidev5R36;
  logic [0:0] callResR136;
  logic [106:0] gzdLLziMainzidev5R37;
  logic [0:0] callResR137;
  logic [106:0] gzdLLziMainzidev5R38;
  logic [0:0] callResR138;
  logic [106:0] gzdLLziMainzidev5R39;
  logic [0:0] callResR139;
  logic [106:0] gzdLLziMainzidev5R40;
  logic [0:0] callResR140;
  logic [106:0] gzdLLziMainzidev5R41;
  logic [0:0] callResR141;
  logic [106:0] gzdLLziMainzidev5R42;
  logic [0:0] callResR142;
  logic [106:0] gzdLLziMainzidev5R43;
  logic [0:0] callResR143;
  logic [106:0] gzdLLziMainzidev5R44;
  logic [0:0] callResR144;
  logic [106:0] gzdLLziMainzidev5R45;
  logic [0:0] callResR145;
  logic [106:0] gzdLLziMainzidev5R46;
  logic [0:0] callResR146;
  logic [106:0] gzdLLziMainzidev5R47;
  logic [0:0] callResR147;
  logic [106:0] gzdLLziMainzidev5R48;
  logic [0:0] callResR148;
  logic [106:0] gzdLLziMainzidev5R49;
  logic [0:0] callResR149;
  logic [106:0] gzdLLziMainzidev5R50;
  logic [0:0] callResR150;
  logic [106:0] gzdLLziMainzidev5R51;
  logic [0:0] callResR151;
  logic [106:0] gzdLLziMainzidev5R52;
  logic [0:0] callResR152;
  logic [106:0] gzdLLziMainzidev5R53;
  logic [0:0] callResR153;
  logic [106:0] gzdLLziMainzidev5R54;
  logic [0:0] callResR154;
  logic [106:0] gzdLLziMainzidev5R55;
  logic [0:0] callResR155;
  logic [106:0] gzdLLziMainzidev5R56;
  logic [0:0] callResR156;
  logic [106:0] gzdLLziMainzidev5R57;
  logic [0:0] callResR157;
  logic [106:0] gzdLLziMainzidev5R58;
  logic [0:0] callResR158;
  logic [106:0] gzdLLziMainzidev5R59;
  logic [0:0] callResR159;
  logic [106:0] gzdLLziMainzidev5R60;
  logic [0:0] callResR160;
  logic [106:0] gzdLLziMainzidev5R61;
  logic [0:0] callResR161;
  logic [106:0] gzdLLziMainzidev5R62;
  logic [0:0] callResR162;
  logic [106:0] gzdLLziMainzidev5R63;
  logic [0:0] callResR163;
  logic [106:0] gzdLLziMainzidev5R64;
  logic [0:0] callResR164;
  logic [106:0] gzdLLziMainzidev5R65;
  logic [0:0] callResR165;
  logic [106:0] gzdLLziMainzidev5R66;
  logic [0:0] callResR166;
  logic [106:0] gzdLLziMainzidev5R67;
  logic [0:0] callResR167;
  logic [106:0] gzdLLziMainzidev5R68;
  logic [0:0] callResR168;
  logic [106:0] gzdLLziMainzidev5R69;
  logic [0:0] callResR169;
  logic [106:0] gzdLLziMainzidev5R70;
  logic [0:0] callResR170;
  logic [106:0] gzdLLziMainzidev5R71;
  logic [0:0] callResR171;
  logic [106:0] gzdLLziMainzidev5R72;
  logic [0:0] callResR172;
  logic [106:0] gzdLLziMainzidev5R73;
  logic [0:0] callResR173;
  logic [106:0] gzdLLziMainzidev5R74;
  logic [0:0] callResR174;
  logic [106:0] gzdLLziMainzidev5R75;
  logic [0:0] callResR175;
  logic [106:0] gzdLLziMainzidev5R76;
  logic [0:0] callResR176;
  logic [106:0] gzdLLziMainzidev5R77;
  logic [0:0] callResR177;
  logic [106:0] gzdLLziMainzidev5R78;
  logic [0:0] callResR178;
  logic [106:0] gzdLLziMainzidev5R79;
  logic [0:0] callResR179;
  logic [106:0] gzdLLziMainzidev5R80;
  logic [0:0] callResR180;
  logic [106:0] gzdLLziMainzidev5R81;
  logic [0:0] callResR181;
  logic [106:0] gzdLLziMainzidev5R82;
  logic [0:0] callResR182;
  logic [106:0] gzdLLziMainzidev5R83;
  logic [0:0] callResR183;
  logic [106:0] gzdLLziMainzidev5R84;
  logic [0:0] callResR184;
  logic [106:0] gzdLLziMainzidev5R85;
  logic [0:0] callResR185;
  logic [106:0] gzdLLziMainzidev5R86;
  logic [0:0] callResR186;
  logic [106:0] gzdLLziMainzidev5R87;
  logic [0:0] callResR187;
  logic [106:0] gzdLLziMainzidev5R88;
  logic [0:0] callResR188;
  logic [106:0] gzdLLziMainzidev5R89;
  logic [0:0] callResR189;
  logic [106:0] gzdLLziMainzidev5R90;
  logic [0:0] callResR190;
  logic [106:0] gzdLLziMainzidev5R91;
  logic [0:0] callResR191;
  logic [106:0] gzdLLziMainzidev5R92;
  logic [0:0] callResR192;
  logic [106:0] gzdLLziMainzidev5R93;
  logic [0:0] callResR193;
  logic [106:0] gzdLLziMainzidev5R94;
  logic [0:0] callResR194;
  logic [106:0] gzdLLziMainzidev5R95;
  logic [0:0] callResR195;
  logic [106:0] gzdLLziMainzidev5R96;
  logic [0:0] callResR196;
  logic [106:0] gzdLLziMainzidev5R97;
  logic [0:0] callResR197;
  logic [106:0] gzdLLziMainzidev5R98;
  logic [0:0] callResR198;
  logic [106:0] gzdLLziMainzidev5R99;
  logic [0:0] callResR199;
  logic [106:0] gzdLLziMainzidev8;
  logic [0:0] callResR200;
  logic [106:0] gzdLLziMainzidev8R1;
  logic [0:0] callResR201;
  logic [106:0] gzdLLziMainzidev8R2;
  logic [0:0] callResR202;
  logic [106:0] gzdLLziMainzidev8R3;
  logic [0:0] callResR203;
  logic [106:0] gzdLLziMainzidev8R4;
  logic [0:0] callResR204;
  logic [106:0] gzdLLziMainzidev8R5;
  logic [0:0] callResR205;
  logic [106:0] gzdLLziMainzidev8R6;
  logic [0:0] callResR206;
  logic [106:0] gzdLLziMainzidev8R7;
  logic [0:0] callResR207;
  logic [106:0] gzdLLziMainzidev8R8;
  logic [0:0] callResR208;
  logic [106:0] gzdLLziMainzidev8R9;
  logic [0:0] callResR209;
  logic [106:0] gzdLLziMainzidev8R10;
  logic [0:0] callResR210;
  logic [106:0] gzdLLziMainzidev8R11;
  logic [0:0] callResR211;
  logic [106:0] gzdLLziMainzidev8R12;
  logic [0:0] callResR212;
  logic [106:0] gzdLLziMainzidev8R13;
  logic [0:0] callResR213;
  logic [106:0] gzdLLziMainzidev8R14;
  logic [0:0] callResR214;
  logic [106:0] gzdLLziMainzidev8R15;
  logic [0:0] callResR215;
  logic [106:0] gzdLLziMainzidev8R16;
  logic [0:0] callResR216;
  logic [106:0] gzdLLziMainzidev8R17;
  logic [0:0] callResR217;
  logic [106:0] gzdLLziMainzidev8R18;
  logic [0:0] callResR218;
  logic [106:0] gzdLLziMainzidev8R19;
  logic [0:0] callResR219;
  logic [106:0] gzdLLziMainzidev8R20;
  logic [0:0] callResR220;
  logic [106:0] gzdLLziMainzidev8R21;
  logic [0:0] callResR221;
  logic [106:0] gzdLLziMainzidev8R22;
  logic [0:0] callResR222;
  logic [106:0] gzdLLziMainzidev8R23;
  logic [0:0] callResR223;
  logic [106:0] gzdLLziMainzidev8R24;
  logic [0:0] callResR224;
  logic [106:0] gzdLLziMainzidev8R25;
  logic [0:0] callResR225;
  logic [106:0] gzdLLziMainzidev8R26;
  logic [0:0] callResR226;
  logic [106:0] gzdLLziMainzidev8R27;
  logic [0:0] callResR227;
  logic [106:0] gzdLLziMainzidev8R28;
  logic [0:0] callResR228;
  logic [106:0] gzdLLziMainzidev8R29;
  logic [0:0] callResR229;
  logic [106:0] gzdLLziMainzidev8R30;
  logic [0:0] callResR230;
  logic [106:0] gzdLLziMainzidev8R31;
  logic [0:0] callResR231;
  logic [106:0] gzdLLziMainzidev8R32;
  logic [0:0] callResR232;
  logic [106:0] gzdLLziMainzidev8R33;
  logic [0:0] callResR233;
  logic [106:0] gzdLLziMainzidev8R34;
  logic [0:0] callResR234;
  logic [106:0] gzdLLziMainzidev8R35;
  logic [0:0] callResR235;
  logic [106:0] gzdLLziMainzidev8R36;
  logic [0:0] callResR236;
  logic [106:0] gzdLLziMainzidev8R37;
  logic [0:0] callResR237;
  logic [106:0] gzdLLziMainzidev8R38;
  logic [0:0] callResR238;
  logic [106:0] gzdLLziMainzidev8R39;
  logic [0:0] callResR239;
  logic [106:0] gzdLLziMainzidev8R40;
  logic [0:0] callResR240;
  logic [106:0] gzdLLziMainzidev8R41;
  logic [0:0] callResR241;
  logic [106:0] gzdLLziMainzidev8R42;
  logic [0:0] callResR242;
  logic [106:0] gzdLLziMainzidev8R43;
  logic [0:0] callResR243;
  logic [106:0] gzdLLziMainzidev8R44;
  logic [0:0] callResR244;
  logic [106:0] gzdLLziMainzidev8R45;
  logic [0:0] callResR245;
  logic [106:0] gzdLLziMainzidev8R46;
  logic [0:0] callResR246;
  logic [106:0] gzdLLziMainzidev8R47;
  logic [0:0] callResR247;
  logic [106:0] gzdLLziMainzidev8R48;
  logic [0:0] callResR248;
  logic [106:0] gzdLLziMainzidev8R49;
  logic [0:0] callResR249;
  logic [106:0] gzdLLziMainzidev8R50;
  logic [0:0] callResR250;
  logic [106:0] gzdLLziMainzidev8R51;
  logic [0:0] callResR251;
  logic [106:0] gzdLLziMainzidev8R52;
  logic [0:0] callResR252;
  logic [106:0] gzdLLziMainzidev8R53;
  logic [0:0] callResR253;
  logic [106:0] gzdLLziMainzidev8R54;
  logic [0:0] callResR254;
  logic [106:0] gzdLLziMainzidev8R55;
  logic [0:0] callResR255;
  logic [106:0] gzdLLziMainzidev8R56;
  logic [0:0] callResR256;
  logic [106:0] gzdLLziMainzidev8R57;
  logic [0:0] callResR257;
  logic [106:0] gzdLLziMainzidev8R58;
  logic [0:0] callResR258;
  logic [106:0] gzdLLziMainzidev8R59;
  logic [0:0] callResR259;
  logic [106:0] gzdLLziMainzidev8R60;
  logic [0:0] callResR260;
  logic [106:0] gzdLLziMainzidev8R61;
  logic [0:0] callResR261;
  logic [106:0] gzdLLziMainzidev8R62;
  logic [0:0] callResR262;
  logic [106:0] gzdLLziMainzidev8R63;
  logic [0:0] callResR263;
  logic [106:0] gzdLLziMainzidev8R64;
  logic [0:0] callResR264;
  logic [106:0] gzdLLziMainzidev8R65;
  logic [0:0] callResR265;
  logic [106:0] gzdLLziMainzidev8R66;
  logic [0:0] callResR266;
  logic [106:0] gzdLLziMainzidev8R67;
  logic [0:0] callResR267;
  logic [106:0] gzdLLziMainzidev8R68;
  logic [0:0] callResR268;
  logic [106:0] gzdLLziMainzidev8R69;
  logic [0:0] callResR269;
  logic [106:0] gzdLLziMainzidev8R70;
  logic [0:0] callResR270;
  logic [106:0] gzdLLziMainzidev8R71;
  logic [0:0] callResR271;
  logic [106:0] gzdLLziMainzidev8R72;
  logic [0:0] callResR272;
  logic [106:0] gzdLLziMainzidev8R73;
  logic [0:0] callResR273;
  logic [106:0] gzdLLziMainzidev8R74;
  logic [0:0] callResR274;
  logic [106:0] gzdLLziMainzidev8R75;
  logic [0:0] callResR275;
  logic [106:0] gzdLLziMainzidev8R76;
  logic [0:0] callResR276;
  logic [106:0] gzdLLziMainzidev8R77;
  logic [0:0] callResR277;
  logic [106:0] gzdLLziMainzidev8R78;
  logic [0:0] callResR278;
  logic [106:0] gzdLLziMainzidev8R79;
  logic [0:0] callResR279;
  logic [106:0] gzdLLziMainzidev8R80;
  logic [0:0] callResR280;
  logic [106:0] gzdLLziMainzidev8R81;
  logic [0:0] callResR281;
  logic [106:0] gzdLLziMainzidev8R82;
  logic [0:0] callResR282;
  logic [106:0] gzdLLziMainzidev8R83;
  logic [0:0] callResR283;
  logic [106:0] gzdLLziMainzidev8R84;
  logic [0:0] callResR284;
  logic [106:0] gzdLLziMainzidev8R85;
  logic [0:0] callResR285;
  logic [106:0] gzdLLziMainzidev8R86;
  logic [0:0] callResR286;
  logic [106:0] gzdLLziMainzidev8R87;
  logic [0:0] callResR287;
  logic [106:0] gzdLLziMainzidev8R88;
  logic [0:0] callResR288;
  logic [106:0] gzdLLziMainzidev8R89;
  logic [0:0] callResR289;
  logic [106:0] gzdLLziMainzidev8R90;
  logic [0:0] callResR290;
  logic [106:0] gzdLLziMainzidev8R91;
  logic [0:0] callResR291;
  logic [106:0] gzdLLziMainzidev8R92;
  logic [0:0] callResR292;
  logic [106:0] gzdLLziMainzidev8R93;
  logic [0:0] callResR293;
  logic [106:0] gzdLLziMainzidev8R94;
  logic [0:0] callResR294;
  logic [106:0] gzdLLziMainzidev8R95;
  logic [0:0] callResR295;
  logic [106:0] gzdLLziMainzidev8R96;
  logic [0:0] callResR296;
  logic [106:0] gzdLLziMainzidev8R97;
  logic [0:0] callResR297;
  logic [106:0] gzdLLziMainzidev8R98;
  logic [0:0] callResR298;
  logic [106:0] gzdLLziMainzidev8R99;
  logic [0:0] callResR299;
  logic [106:0] gzdLLziMainzidev11;
  logic [0:0] callResR300;
  logic [106:0] gzdLLziMainzidev11R1;
  logic [0:0] callResR301;
  logic [106:0] gzdLLziMainzidev11R2;
  logic [0:0] callResR302;
  logic [106:0] gzdLLziMainzidev11R3;
  logic [0:0] callResR303;
  logic [106:0] gzdLLziMainzidev11R4;
  logic [0:0] callResR304;
  logic [106:0] gzdLLziMainzidev11R5;
  logic [0:0] callResR305;
  logic [106:0] gzdLLziMainzidev11R6;
  logic [0:0] callResR306;
  logic [106:0] gzdLLziMainzidev11R7;
  logic [0:0] callResR307;
  logic [106:0] gzdLLziMainzidev11R8;
  logic [0:0] callResR308;
  logic [106:0] gzdLLziMainzidev11R9;
  logic [0:0] callResR309;
  logic [106:0] gzdLLziMainzidev11R10;
  logic [0:0] callResR310;
  logic [106:0] gzdLLziMainzidev11R11;
  logic [0:0] callResR311;
  logic [106:0] gzdLLziMainzidev11R12;
  logic [0:0] callResR312;
  logic [106:0] gzdLLziMainzidev11R13;
  logic [0:0] callResR313;
  logic [106:0] gzdLLziMainzidev11R14;
  logic [0:0] callResR314;
  logic [106:0] gzdLLziMainzidev11R15;
  logic [0:0] callResR315;
  logic [106:0] gzdLLziMainzidev11R16;
  logic [0:0] callResR316;
  logic [106:0] gzdLLziMainzidev11R17;
  logic [0:0] callResR317;
  logic [106:0] gzdLLziMainzidev11R18;
  logic [0:0] callResR318;
  logic [106:0] gzdLLziMainzidev11R19;
  logic [0:0] callResR319;
  logic [106:0] gzdLLziMainzidev11R20;
  logic [0:0] callResR320;
  logic [106:0] gzdLLziMainzidev11R21;
  logic [0:0] callResR321;
  logic [106:0] gzdLLziMainzidev11R22;
  logic [0:0] callResR322;
  logic [106:0] gzdLLziMainzidev11R23;
  logic [0:0] callResR323;
  logic [106:0] gzdLLziMainzidev11R24;
  logic [0:0] callResR324;
  logic [106:0] gzdLLziMainzidev11R25;
  logic [0:0] callResR325;
  logic [106:0] gzdLLziMainzidev11R26;
  logic [0:0] callResR326;
  logic [106:0] gzdLLziMainzidev11R27;
  logic [0:0] callResR327;
  logic [106:0] gzdLLziMainzidev11R28;
  logic [0:0] callResR328;
  logic [106:0] gzdLLziMainzidev11R29;
  logic [0:0] callResR329;
  logic [106:0] gzdLLziMainzidev11R30;
  logic [0:0] callResR330;
  logic [106:0] gzdLLziMainzidev11R31;
  logic [0:0] callResR331;
  logic [106:0] gzdLLziMainzidev11R32;
  logic [0:0] callResR332;
  logic [106:0] gzdLLziMainzidev11R33;
  logic [0:0] callResR333;
  logic [106:0] gzdLLziMainzidev11R34;
  logic [0:0] callResR334;
  logic [106:0] gzdLLziMainzidev11R35;
  logic [0:0] callResR335;
  logic [106:0] gzdLLziMainzidev11R36;
  logic [0:0] callResR336;
  logic [106:0] gzdLLziMainzidev11R37;
  logic [0:0] callResR337;
  logic [106:0] gzdLLziMainzidev11R38;
  logic [0:0] callResR338;
  logic [106:0] gzdLLziMainzidev11R39;
  logic [0:0] callResR339;
  logic [106:0] gzdLLziMainzidev11R40;
  logic [0:0] callResR340;
  logic [106:0] gzdLLziMainzidev11R41;
  logic [0:0] callResR341;
  logic [106:0] gzdLLziMainzidev11R42;
  logic [0:0] callResR342;
  logic [106:0] gzdLLziMainzidev11R43;
  logic [0:0] callResR343;
  logic [106:0] gzdLLziMainzidev11R44;
  logic [0:0] callResR344;
  logic [106:0] gzdLLziMainzidev11R45;
  logic [0:0] callResR345;
  logic [106:0] gzdLLziMainzidev11R46;
  logic [0:0] callResR346;
  logic [106:0] gzdLLziMainzidev11R47;
  logic [0:0] callResR347;
  logic [106:0] gzdLLziMainzidev11R48;
  logic [0:0] callResR348;
  logic [106:0] gzdLLziMainzidev11R49;
  logic [0:0] callResR349;
  logic [106:0] gzdLLziMainzidev11R50;
  logic [0:0] callResR350;
  logic [106:0] gzdLLziMainzidev11R51;
  logic [0:0] callResR351;
  logic [106:0] gzdLLziMainzidev11R52;
  logic [0:0] callResR352;
  logic [106:0] gzdLLziMainzidev11R53;
  logic [0:0] callResR353;
  logic [106:0] gzdLLziMainzidev11R54;
  logic [0:0] callResR354;
  logic [106:0] gzdLLziMainzidev11R55;
  logic [0:0] callResR355;
  logic [106:0] gzdLLziMainzidev11R56;
  logic [0:0] callResR356;
  logic [106:0] gzdLLziMainzidev11R57;
  logic [0:0] callResR357;
  logic [106:0] gzdLLziMainzidev11R58;
  logic [0:0] callResR358;
  logic [106:0] gzdLLziMainzidev11R59;
  logic [0:0] callResR359;
  logic [106:0] gzdLLziMainzidev11R60;
  logic [0:0] callResR360;
  logic [106:0] gzdLLziMainzidev11R61;
  logic [0:0] callResR361;
  logic [106:0] gzdLLziMainzidev11R62;
  logic [0:0] callResR362;
  logic [106:0] gzdLLziMainzidev11R63;
  logic [0:0] callResR363;
  logic [106:0] gzdLLziMainzidev11R64;
  logic [0:0] callResR364;
  logic [106:0] gzdLLziMainzidev11R65;
  logic [0:0] callResR365;
  logic [106:0] gzdLLziMainzidev11R66;
  logic [0:0] callResR366;
  logic [106:0] gzdLLziMainzidev11R67;
  logic [0:0] callResR367;
  logic [106:0] gzdLLziMainzidev11R68;
  logic [0:0] callResR368;
  logic [106:0] gzdLLziMainzidev11R69;
  logic [0:0] callResR369;
  logic [106:0] gzdLLziMainzidev11R70;
  logic [0:0] callResR370;
  logic [106:0] gzdLLziMainzidev11R71;
  logic [0:0] callResR371;
  logic [106:0] gzdLLziMainzidev11R72;
  logic [0:0] callResR372;
  logic [106:0] gzdLLziMainzidev11R73;
  logic [0:0] callResR373;
  logic [106:0] gzdLLziMainzidev11R74;
  logic [0:0] callResR374;
  logic [106:0] gzdLLziMainzidev11R75;
  logic [0:0] callResR375;
  logic [106:0] gzdLLziMainzidev11R76;
  logic [0:0] callResR376;
  logic [106:0] gzdLLziMainzidev11R77;
  logic [0:0] callResR377;
  logic [106:0] gzdLLziMainzidev11R78;
  logic [0:0] callResR378;
  logic [106:0] gzdLLziMainzidev11R79;
  logic [0:0] callResR379;
  logic [106:0] gzdLLziMainzidev11R80;
  logic [0:0] callResR380;
  logic [106:0] gzdLLziMainzidev11R81;
  logic [0:0] callResR381;
  logic [106:0] gzdLLziMainzidev11R82;
  logic [0:0] callResR382;
  logic [106:0] gzdLLziMainzidev11R83;
  logic [0:0] callResR383;
  logic [106:0] gzdLLziMainzidev11R84;
  logic [0:0] callResR384;
  logic [106:0] gzdLLziMainzidev11R85;
  logic [0:0] callResR385;
  logic [106:0] gzdLLziMainzidev11R86;
  logic [0:0] callResR386;
  logic [106:0] gzdLLziMainzidev11R87;
  logic [0:0] callResR387;
  logic [106:0] gzdLLziMainzidev11R88;
  logic [0:0] callResR388;
  logic [106:0] gzdLLziMainzidev11R89;
  logic [0:0] callResR389;
  logic [106:0] gzdLLziMainzidev11R90;
  logic [0:0] callResR390;
  logic [106:0] gzdLLziMainzidev11R91;
  logic [0:0] callResR391;
  logic [106:0] gzdLLziMainzidev11R92;
  logic [0:0] callResR392;
  logic [106:0] gzdLLziMainzidev11R93;
  logic [0:0] callResR393;
  logic [106:0] gzdLLziMainzidev11R94;
  logic [0:0] callResR394;
  logic [106:0] gzdLLziMainzidev11R95;
  logic [0:0] callResR395;
  logic [106:0] gzdLLziMainzidev11R96;
  logic [0:0] callResR396;
  logic [106:0] gzdLLziMainzidev11R97;
  logic [0:0] callResR397;
  logic [106:0] gzdLLziMainzidev11R98;
  logic [0:0] callResR398;
  logic [106:0] gzdLLziMainzidev11R99;
  logic [0:0] callResR399;
  logic [0:0] __continue;
  logic [99:0] __resumption_tag;
  logic [99:0] __resumption_tag_next;
  assign gMainzidev = __resumption_tag;
  assign gzdLLziMainzidev2 = {gMainzidev[99:0], 7'h00};
  zdLLziMainzidev2  zdLLziMainzidev2 (gzdLLziMainzidev2[106:7], gzdLLziMainzidev2[6:0], callRes);
  assign gzdLLziMainzidev2R1 = {gMainzidev[99:0], 7'h01};
  zdLLziMainzidev2  zdLLziMainzidev2R1 (gzdLLziMainzidev2R1[106:7], gzdLLziMainzidev2R1[6:0], callResR1);
  assign gzdLLziMainzidev2R2 = {gMainzidev[99:0], 7'h02};
  zdLLziMainzidev2  zdLLziMainzidev2R2 (gzdLLziMainzidev2R2[106:7], gzdLLziMainzidev2R2[6:0], callResR2);
  assign gzdLLziMainzidev2R3 = {gMainzidev[99:0], 7'h03};
  zdLLziMainzidev2  zdLLziMainzidev2R3 (gzdLLziMainzidev2R3[106:7], gzdLLziMainzidev2R3[6:0], callResR3);
  assign gzdLLziMainzidev2R4 = {gMainzidev[99:0], 7'h04};
  zdLLziMainzidev2  zdLLziMainzidev2R4 (gzdLLziMainzidev2R4[106:7], gzdLLziMainzidev2R4[6:0], callResR4);
  assign gzdLLziMainzidev2R5 = {gMainzidev[99:0], 7'h05};
  zdLLziMainzidev2  zdLLziMainzidev2R5 (gzdLLziMainzidev2R5[106:7], gzdLLziMainzidev2R5[6:0], callResR5);
  assign gzdLLziMainzidev2R6 = {gMainzidev[99:0], 7'h06};
  zdLLziMainzidev2  zdLLziMainzidev2R6 (gzdLLziMainzidev2R6[106:7], gzdLLziMainzidev2R6[6:0], callResR6);
  assign gzdLLziMainzidev2R7 = {gMainzidev[99:0], 7'h07};
  zdLLziMainzidev2  zdLLziMainzidev2R7 (gzdLLziMainzidev2R7[106:7], gzdLLziMainzidev2R7[6:0], callResR7);
  assign gzdLLziMainzidev2R8 = {gMainzidev[99:0], 7'h08};
  zdLLziMainzidev2  zdLLziMainzidev2R8 (gzdLLziMainzidev2R8[106:7], gzdLLziMainzidev2R8[6:0], callResR8);
  assign gzdLLziMainzidev2R9 = {gMainzidev[99:0], 7'h09};
  zdLLziMainzidev2  zdLLziMainzidev2R9 (gzdLLziMainzidev2R9[106:7], gzdLLziMainzidev2R9[6:0], callResR9);
  assign gzdLLziMainzidev2R10 = {gMainzidev[99:0], 7'h0a};
  zdLLziMainzidev2  zdLLziMainzidev2R10 (gzdLLziMainzidev2R10[106:7], gzdLLziMainzidev2R10[6:0], callResR10);
  assign gzdLLziMainzidev2R11 = {gMainzidev[99:0], 7'h0b};
  zdLLziMainzidev2  zdLLziMainzidev2R11 (gzdLLziMainzidev2R11[106:7], gzdLLziMainzidev2R11[6:0], callResR11);
  assign gzdLLziMainzidev2R12 = {gMainzidev[99:0], 7'h0c};
  zdLLziMainzidev2  zdLLziMainzidev2R12 (gzdLLziMainzidev2R12[106:7], gzdLLziMainzidev2R12[6:0], callResR12);
  assign gzdLLziMainzidev2R13 = {gMainzidev[99:0], 7'h0d};
  zdLLziMainzidev2  zdLLziMainzidev2R13 (gzdLLziMainzidev2R13[106:7], gzdLLziMainzidev2R13[6:0], callResR13);
  assign gzdLLziMainzidev2R14 = {gMainzidev[99:0], 7'h0e};
  zdLLziMainzidev2  zdLLziMainzidev2R14 (gzdLLziMainzidev2R14[106:7], gzdLLziMainzidev2R14[6:0], callResR14);
  assign gzdLLziMainzidev2R15 = {gMainzidev[99:0], 7'h0f};
  zdLLziMainzidev2  zdLLziMainzidev2R15 (gzdLLziMainzidev2R15[106:7], gzdLLziMainzidev2R15[6:0], callResR15);
  assign gzdLLziMainzidev2R16 = {gMainzidev[99:0], 7'h10};
  zdLLziMainzidev2  zdLLziMainzidev2R16 (gzdLLziMainzidev2R16[106:7], gzdLLziMainzidev2R16[6:0], callResR16);
  assign gzdLLziMainzidev2R17 = {gMainzidev[99:0], 7'h11};
  zdLLziMainzidev2  zdLLziMainzidev2R17 (gzdLLziMainzidev2R17[106:7], gzdLLziMainzidev2R17[6:0], callResR17);
  assign gzdLLziMainzidev2R18 = {gMainzidev[99:0], 7'h12};
  zdLLziMainzidev2  zdLLziMainzidev2R18 (gzdLLziMainzidev2R18[106:7], gzdLLziMainzidev2R18[6:0], callResR18);
  assign gzdLLziMainzidev2R19 = {gMainzidev[99:0], 7'h13};
  zdLLziMainzidev2  zdLLziMainzidev2R19 (gzdLLziMainzidev2R19[106:7], gzdLLziMainzidev2R19[6:0], callResR19);
  assign gzdLLziMainzidev2R20 = {gMainzidev[99:0], 7'h14};
  zdLLziMainzidev2  zdLLziMainzidev2R20 (gzdLLziMainzidev2R20[106:7], gzdLLziMainzidev2R20[6:0], callResR20);
  assign gzdLLziMainzidev2R21 = {gMainzidev[99:0], 7'h15};
  zdLLziMainzidev2  zdLLziMainzidev2R21 (gzdLLziMainzidev2R21[106:7], gzdLLziMainzidev2R21[6:0], callResR21);
  assign gzdLLziMainzidev2R22 = {gMainzidev[99:0], 7'h16};
  zdLLziMainzidev2  zdLLziMainzidev2R22 (gzdLLziMainzidev2R22[106:7], gzdLLziMainzidev2R22[6:0], callResR22);
  assign gzdLLziMainzidev2R23 = {gMainzidev[99:0], 7'h17};
  zdLLziMainzidev2  zdLLziMainzidev2R23 (gzdLLziMainzidev2R23[106:7], gzdLLziMainzidev2R23[6:0], callResR23);
  assign gzdLLziMainzidev2R24 = {gMainzidev[99:0], 7'h18};
  zdLLziMainzidev2  zdLLziMainzidev2R24 (gzdLLziMainzidev2R24[106:7], gzdLLziMainzidev2R24[6:0], callResR24);
  assign gzdLLziMainzidev2R25 = {gMainzidev[99:0], 7'h19};
  zdLLziMainzidev2  zdLLziMainzidev2R25 (gzdLLziMainzidev2R25[106:7], gzdLLziMainzidev2R25[6:0], callResR25);
  assign gzdLLziMainzidev2R26 = {gMainzidev[99:0], 7'h1a};
  zdLLziMainzidev2  zdLLziMainzidev2R26 (gzdLLziMainzidev2R26[106:7], gzdLLziMainzidev2R26[6:0], callResR26);
  assign gzdLLziMainzidev2R27 = {gMainzidev[99:0], 7'h1b};
  zdLLziMainzidev2  zdLLziMainzidev2R27 (gzdLLziMainzidev2R27[106:7], gzdLLziMainzidev2R27[6:0], callResR27);
  assign gzdLLziMainzidev2R28 = {gMainzidev[99:0], 7'h1c};
  zdLLziMainzidev2  zdLLziMainzidev2R28 (gzdLLziMainzidev2R28[106:7], gzdLLziMainzidev2R28[6:0], callResR28);
  assign gzdLLziMainzidev2R29 = {gMainzidev[99:0], 7'h1d};
  zdLLziMainzidev2  zdLLziMainzidev2R29 (gzdLLziMainzidev2R29[106:7], gzdLLziMainzidev2R29[6:0], callResR29);
  assign gzdLLziMainzidev2R30 = {gMainzidev[99:0], 7'h1e};
  zdLLziMainzidev2  zdLLziMainzidev2R30 (gzdLLziMainzidev2R30[106:7], gzdLLziMainzidev2R30[6:0], callResR30);
  assign gzdLLziMainzidev2R31 = {gMainzidev[99:0], 7'h1f};
  zdLLziMainzidev2  zdLLziMainzidev2R31 (gzdLLziMainzidev2R31[106:7], gzdLLziMainzidev2R31[6:0], callResR31);
  assign gzdLLziMainzidev2R32 = {gMainzidev[99:0], 7'h20};
  zdLLziMainzidev2  zdLLziMainzidev2R32 (gzdLLziMainzidev2R32[106:7], gzdLLziMainzidev2R32[6:0], callResR32);
  assign gzdLLziMainzidev2R33 = {gMainzidev[99:0], 7'h21};
  zdLLziMainzidev2  zdLLziMainzidev2R33 (gzdLLziMainzidev2R33[106:7], gzdLLziMainzidev2R33[6:0], callResR33);
  assign gzdLLziMainzidev2R34 = {gMainzidev[99:0], 7'h22};
  zdLLziMainzidev2  zdLLziMainzidev2R34 (gzdLLziMainzidev2R34[106:7], gzdLLziMainzidev2R34[6:0], callResR34);
  assign gzdLLziMainzidev2R35 = {gMainzidev[99:0], 7'h23};
  zdLLziMainzidev2  zdLLziMainzidev2R35 (gzdLLziMainzidev2R35[106:7], gzdLLziMainzidev2R35[6:0], callResR35);
  assign gzdLLziMainzidev2R36 = {gMainzidev[99:0], 7'h24};
  zdLLziMainzidev2  zdLLziMainzidev2R36 (gzdLLziMainzidev2R36[106:7], gzdLLziMainzidev2R36[6:0], callResR36);
  assign gzdLLziMainzidev2R37 = {gMainzidev[99:0], 7'h25};
  zdLLziMainzidev2  zdLLziMainzidev2R37 (gzdLLziMainzidev2R37[106:7], gzdLLziMainzidev2R37[6:0], callResR37);
  assign gzdLLziMainzidev2R38 = {gMainzidev[99:0], 7'h26};
  zdLLziMainzidev2  zdLLziMainzidev2R38 (gzdLLziMainzidev2R38[106:7], gzdLLziMainzidev2R38[6:0], callResR38);
  assign gzdLLziMainzidev2R39 = {gMainzidev[99:0], 7'h27};
  zdLLziMainzidev2  zdLLziMainzidev2R39 (gzdLLziMainzidev2R39[106:7], gzdLLziMainzidev2R39[6:0], callResR39);
  assign gzdLLziMainzidev2R40 = {gMainzidev[99:0], 7'h28};
  zdLLziMainzidev2  zdLLziMainzidev2R40 (gzdLLziMainzidev2R40[106:7], gzdLLziMainzidev2R40[6:0], callResR40);
  assign gzdLLziMainzidev2R41 = {gMainzidev[99:0], 7'h29};
  zdLLziMainzidev2  zdLLziMainzidev2R41 (gzdLLziMainzidev2R41[106:7], gzdLLziMainzidev2R41[6:0], callResR41);
  assign gzdLLziMainzidev2R42 = {gMainzidev[99:0], 7'h2a};
  zdLLziMainzidev2  zdLLziMainzidev2R42 (gzdLLziMainzidev2R42[106:7], gzdLLziMainzidev2R42[6:0], callResR42);
  assign gzdLLziMainzidev2R43 = {gMainzidev[99:0], 7'h2b};
  zdLLziMainzidev2  zdLLziMainzidev2R43 (gzdLLziMainzidev2R43[106:7], gzdLLziMainzidev2R43[6:0], callResR43);
  assign gzdLLziMainzidev2R44 = {gMainzidev[99:0], 7'h2c};
  zdLLziMainzidev2  zdLLziMainzidev2R44 (gzdLLziMainzidev2R44[106:7], gzdLLziMainzidev2R44[6:0], callResR44);
  assign gzdLLziMainzidev2R45 = {gMainzidev[99:0], 7'h2d};
  zdLLziMainzidev2  zdLLziMainzidev2R45 (gzdLLziMainzidev2R45[106:7], gzdLLziMainzidev2R45[6:0], callResR45);
  assign gzdLLziMainzidev2R46 = {gMainzidev[99:0], 7'h2e};
  zdLLziMainzidev2  zdLLziMainzidev2R46 (gzdLLziMainzidev2R46[106:7], gzdLLziMainzidev2R46[6:0], callResR46);
  assign gzdLLziMainzidev2R47 = {gMainzidev[99:0], 7'h2f};
  zdLLziMainzidev2  zdLLziMainzidev2R47 (gzdLLziMainzidev2R47[106:7], gzdLLziMainzidev2R47[6:0], callResR47);
  assign gzdLLziMainzidev2R48 = {gMainzidev[99:0], 7'h30};
  zdLLziMainzidev2  zdLLziMainzidev2R48 (gzdLLziMainzidev2R48[106:7], gzdLLziMainzidev2R48[6:0], callResR48);
  assign gzdLLziMainzidev2R49 = {gMainzidev[99:0], 7'h31};
  zdLLziMainzidev2  zdLLziMainzidev2R49 (gzdLLziMainzidev2R49[106:7], gzdLLziMainzidev2R49[6:0], callResR49);
  assign gzdLLziMainzidev2R50 = {gMainzidev[99:0], 7'h32};
  zdLLziMainzidev2  zdLLziMainzidev2R50 (gzdLLziMainzidev2R50[106:7], gzdLLziMainzidev2R50[6:0], callResR50);
  assign gzdLLziMainzidev2R51 = {gMainzidev[99:0], 7'h33};
  zdLLziMainzidev2  zdLLziMainzidev2R51 (gzdLLziMainzidev2R51[106:7], gzdLLziMainzidev2R51[6:0], callResR51);
  assign gzdLLziMainzidev2R52 = {gMainzidev[99:0], 7'h34};
  zdLLziMainzidev2  zdLLziMainzidev2R52 (gzdLLziMainzidev2R52[106:7], gzdLLziMainzidev2R52[6:0], callResR52);
  assign gzdLLziMainzidev2R53 = {gMainzidev[99:0], 7'h35};
  zdLLziMainzidev2  zdLLziMainzidev2R53 (gzdLLziMainzidev2R53[106:7], gzdLLziMainzidev2R53[6:0], callResR53);
  assign gzdLLziMainzidev2R54 = {gMainzidev[99:0], 7'h36};
  zdLLziMainzidev2  zdLLziMainzidev2R54 (gzdLLziMainzidev2R54[106:7], gzdLLziMainzidev2R54[6:0], callResR54);
  assign gzdLLziMainzidev2R55 = {gMainzidev[99:0], 7'h37};
  zdLLziMainzidev2  zdLLziMainzidev2R55 (gzdLLziMainzidev2R55[106:7], gzdLLziMainzidev2R55[6:0], callResR55);
  assign gzdLLziMainzidev2R56 = {gMainzidev[99:0], 7'h38};
  zdLLziMainzidev2  zdLLziMainzidev2R56 (gzdLLziMainzidev2R56[106:7], gzdLLziMainzidev2R56[6:0], callResR56);
  assign gzdLLziMainzidev2R57 = {gMainzidev[99:0], 7'h39};
  zdLLziMainzidev2  zdLLziMainzidev2R57 (gzdLLziMainzidev2R57[106:7], gzdLLziMainzidev2R57[6:0], callResR57);
  assign gzdLLziMainzidev2R58 = {gMainzidev[99:0], 7'h3a};
  zdLLziMainzidev2  zdLLziMainzidev2R58 (gzdLLziMainzidev2R58[106:7], gzdLLziMainzidev2R58[6:0], callResR58);
  assign gzdLLziMainzidev2R59 = {gMainzidev[99:0], 7'h3b};
  zdLLziMainzidev2  zdLLziMainzidev2R59 (gzdLLziMainzidev2R59[106:7], gzdLLziMainzidev2R59[6:0], callResR59);
  assign gzdLLziMainzidev2R60 = {gMainzidev[99:0], 7'h3c};
  zdLLziMainzidev2  zdLLziMainzidev2R60 (gzdLLziMainzidev2R60[106:7], gzdLLziMainzidev2R60[6:0], callResR60);
  assign gzdLLziMainzidev2R61 = {gMainzidev[99:0], 7'h3d};
  zdLLziMainzidev2  zdLLziMainzidev2R61 (gzdLLziMainzidev2R61[106:7], gzdLLziMainzidev2R61[6:0], callResR61);
  assign gzdLLziMainzidev2R62 = {gMainzidev[99:0], 7'h3e};
  zdLLziMainzidev2  zdLLziMainzidev2R62 (gzdLLziMainzidev2R62[106:7], gzdLLziMainzidev2R62[6:0], callResR62);
  assign gzdLLziMainzidev2R63 = {gMainzidev[99:0], 7'h3f};
  zdLLziMainzidev2  zdLLziMainzidev2R63 (gzdLLziMainzidev2R63[106:7], gzdLLziMainzidev2R63[6:0], callResR63);
  assign gzdLLziMainzidev2R64 = {gMainzidev[99:0], 7'h40};
  zdLLziMainzidev2  zdLLziMainzidev2R64 (gzdLLziMainzidev2R64[106:7], gzdLLziMainzidev2R64[6:0], callResR64);
  assign gzdLLziMainzidev2R65 = {gMainzidev[99:0], 7'h41};
  zdLLziMainzidev2  zdLLziMainzidev2R65 (gzdLLziMainzidev2R65[106:7], gzdLLziMainzidev2R65[6:0], callResR65);
  assign gzdLLziMainzidev2R66 = {gMainzidev[99:0], 7'h42};
  zdLLziMainzidev2  zdLLziMainzidev2R66 (gzdLLziMainzidev2R66[106:7], gzdLLziMainzidev2R66[6:0], callResR66);
  assign gzdLLziMainzidev2R67 = {gMainzidev[99:0], 7'h43};
  zdLLziMainzidev2  zdLLziMainzidev2R67 (gzdLLziMainzidev2R67[106:7], gzdLLziMainzidev2R67[6:0], callResR67);
  assign gzdLLziMainzidev2R68 = {gMainzidev[99:0], 7'h44};
  zdLLziMainzidev2  zdLLziMainzidev2R68 (gzdLLziMainzidev2R68[106:7], gzdLLziMainzidev2R68[6:0], callResR68);
  assign gzdLLziMainzidev2R69 = {gMainzidev[99:0], 7'h45};
  zdLLziMainzidev2  zdLLziMainzidev2R69 (gzdLLziMainzidev2R69[106:7], gzdLLziMainzidev2R69[6:0], callResR69);
  assign gzdLLziMainzidev2R70 = {gMainzidev[99:0], 7'h46};
  zdLLziMainzidev2  zdLLziMainzidev2R70 (gzdLLziMainzidev2R70[106:7], gzdLLziMainzidev2R70[6:0], callResR70);
  assign gzdLLziMainzidev2R71 = {gMainzidev[99:0], 7'h47};
  zdLLziMainzidev2  zdLLziMainzidev2R71 (gzdLLziMainzidev2R71[106:7], gzdLLziMainzidev2R71[6:0], callResR71);
  assign gzdLLziMainzidev2R72 = {gMainzidev[99:0], 7'h48};
  zdLLziMainzidev2  zdLLziMainzidev2R72 (gzdLLziMainzidev2R72[106:7], gzdLLziMainzidev2R72[6:0], callResR72);
  assign gzdLLziMainzidev2R73 = {gMainzidev[99:0], 7'h49};
  zdLLziMainzidev2  zdLLziMainzidev2R73 (gzdLLziMainzidev2R73[106:7], gzdLLziMainzidev2R73[6:0], callResR73);
  assign gzdLLziMainzidev2R74 = {gMainzidev[99:0], 7'h4a};
  zdLLziMainzidev2  zdLLziMainzidev2R74 (gzdLLziMainzidev2R74[106:7], gzdLLziMainzidev2R74[6:0], callResR74);
  assign gzdLLziMainzidev2R75 = {gMainzidev[99:0], 7'h4b};
  zdLLziMainzidev2  zdLLziMainzidev2R75 (gzdLLziMainzidev2R75[106:7], gzdLLziMainzidev2R75[6:0], callResR75);
  assign gzdLLziMainzidev2R76 = {gMainzidev[99:0], 7'h4c};
  zdLLziMainzidev2  zdLLziMainzidev2R76 (gzdLLziMainzidev2R76[106:7], gzdLLziMainzidev2R76[6:0], callResR76);
  assign gzdLLziMainzidev2R77 = {gMainzidev[99:0], 7'h4d};
  zdLLziMainzidev2  zdLLziMainzidev2R77 (gzdLLziMainzidev2R77[106:7], gzdLLziMainzidev2R77[6:0], callResR77);
  assign gzdLLziMainzidev2R78 = {gMainzidev[99:0], 7'h4e};
  zdLLziMainzidev2  zdLLziMainzidev2R78 (gzdLLziMainzidev2R78[106:7], gzdLLziMainzidev2R78[6:0], callResR78);
  assign gzdLLziMainzidev2R79 = {gMainzidev[99:0], 7'h4f};
  zdLLziMainzidev2  zdLLziMainzidev2R79 (gzdLLziMainzidev2R79[106:7], gzdLLziMainzidev2R79[6:0], callResR79);
  assign gzdLLziMainzidev2R80 = {gMainzidev[99:0], 7'h50};
  zdLLziMainzidev2  zdLLziMainzidev2R80 (gzdLLziMainzidev2R80[106:7], gzdLLziMainzidev2R80[6:0], callResR80);
  assign gzdLLziMainzidev2R81 = {gMainzidev[99:0], 7'h51};
  zdLLziMainzidev2  zdLLziMainzidev2R81 (gzdLLziMainzidev2R81[106:7], gzdLLziMainzidev2R81[6:0], callResR81);
  assign gzdLLziMainzidev2R82 = {gMainzidev[99:0], 7'h52};
  zdLLziMainzidev2  zdLLziMainzidev2R82 (gzdLLziMainzidev2R82[106:7], gzdLLziMainzidev2R82[6:0], callResR82);
  assign gzdLLziMainzidev2R83 = {gMainzidev[99:0], 7'h53};
  zdLLziMainzidev2  zdLLziMainzidev2R83 (gzdLLziMainzidev2R83[106:7], gzdLLziMainzidev2R83[6:0], callResR83);
  assign gzdLLziMainzidev2R84 = {gMainzidev[99:0], 7'h54};
  zdLLziMainzidev2  zdLLziMainzidev2R84 (gzdLLziMainzidev2R84[106:7], gzdLLziMainzidev2R84[6:0], callResR84);
  assign gzdLLziMainzidev2R85 = {gMainzidev[99:0], 7'h55};
  zdLLziMainzidev2  zdLLziMainzidev2R85 (gzdLLziMainzidev2R85[106:7], gzdLLziMainzidev2R85[6:0], callResR85);
  assign gzdLLziMainzidev2R86 = {gMainzidev[99:0], 7'h56};
  zdLLziMainzidev2  zdLLziMainzidev2R86 (gzdLLziMainzidev2R86[106:7], gzdLLziMainzidev2R86[6:0], callResR86);
  assign gzdLLziMainzidev2R87 = {gMainzidev[99:0], 7'h57};
  zdLLziMainzidev2  zdLLziMainzidev2R87 (gzdLLziMainzidev2R87[106:7], gzdLLziMainzidev2R87[6:0], callResR87);
  assign gzdLLziMainzidev2R88 = {gMainzidev[99:0], 7'h58};
  zdLLziMainzidev2  zdLLziMainzidev2R88 (gzdLLziMainzidev2R88[106:7], gzdLLziMainzidev2R88[6:0], callResR88);
  assign gzdLLziMainzidev2R89 = {gMainzidev[99:0], 7'h59};
  zdLLziMainzidev2  zdLLziMainzidev2R89 (gzdLLziMainzidev2R89[106:7], gzdLLziMainzidev2R89[6:0], callResR89);
  assign gzdLLziMainzidev2R90 = {gMainzidev[99:0], 7'h5a};
  zdLLziMainzidev2  zdLLziMainzidev2R90 (gzdLLziMainzidev2R90[106:7], gzdLLziMainzidev2R90[6:0], callResR90);
  assign gzdLLziMainzidev2R91 = {gMainzidev[99:0], 7'h5b};
  zdLLziMainzidev2  zdLLziMainzidev2R91 (gzdLLziMainzidev2R91[106:7], gzdLLziMainzidev2R91[6:0], callResR91);
  assign gzdLLziMainzidev2R92 = {gMainzidev[99:0], 7'h5c};
  zdLLziMainzidev2  zdLLziMainzidev2R92 (gzdLLziMainzidev2R92[106:7], gzdLLziMainzidev2R92[6:0], callResR92);
  assign gzdLLziMainzidev2R93 = {gMainzidev[99:0], 7'h5d};
  zdLLziMainzidev2  zdLLziMainzidev2R93 (gzdLLziMainzidev2R93[106:7], gzdLLziMainzidev2R93[6:0], callResR93);
  assign gzdLLziMainzidev2R94 = {gMainzidev[99:0], 7'h5e};
  zdLLziMainzidev2  zdLLziMainzidev2R94 (gzdLLziMainzidev2R94[106:7], gzdLLziMainzidev2R94[6:0], callResR94);
  assign gzdLLziMainzidev2R95 = {gMainzidev[99:0], 7'h5f};
  zdLLziMainzidev2  zdLLziMainzidev2R95 (gzdLLziMainzidev2R95[106:7], gzdLLziMainzidev2R95[6:0], callResR95);
  assign gzdLLziMainzidev2R96 = {gMainzidev[99:0], 7'h60};
  zdLLziMainzidev2  zdLLziMainzidev2R96 (gzdLLziMainzidev2R96[106:7], gzdLLziMainzidev2R96[6:0], callResR96);
  assign gzdLLziMainzidev2R97 = {gMainzidev[99:0], 7'h61};
  zdLLziMainzidev2  zdLLziMainzidev2R97 (gzdLLziMainzidev2R97[106:7], gzdLLziMainzidev2R97[6:0], callResR97);
  assign gzdLLziMainzidev2R98 = {gMainzidev[99:0], 7'h62};
  zdLLziMainzidev2  zdLLziMainzidev2R98 (gzdLLziMainzidev2R98[106:7], gzdLLziMainzidev2R98[6:0], callResR98);
  assign gzdLLziMainzidev2R99 = {gMainzidev[99:0], 7'h63};
  zdLLziMainzidev2  zdLLziMainzidev2R99 (gzdLLziMainzidev2R99[106:7], gzdLLziMainzidev2R99[6:0], callResR99);
  assign gzdLLziMainzidev5 = {gMainzidev[99:0], 7'h00};
  zdLLziMainzidev5  zdLLziMainzidev5 (gzdLLziMainzidev5[106:7], gzdLLziMainzidev5[6:0], callResR100);
  assign gzdLLziMainzidev5R1 = {gMainzidev[99:0], 7'h01};
  zdLLziMainzidev5  zdLLziMainzidev5R1 (gzdLLziMainzidev5R1[106:7], gzdLLziMainzidev5R1[6:0], callResR101);
  assign gzdLLziMainzidev5R2 = {gMainzidev[99:0], 7'h02};
  zdLLziMainzidev5  zdLLziMainzidev5R2 (gzdLLziMainzidev5R2[106:7], gzdLLziMainzidev5R2[6:0], callResR102);
  assign gzdLLziMainzidev5R3 = {gMainzidev[99:0], 7'h03};
  zdLLziMainzidev5  zdLLziMainzidev5R3 (gzdLLziMainzidev5R3[106:7], gzdLLziMainzidev5R3[6:0], callResR103);
  assign gzdLLziMainzidev5R4 = {gMainzidev[99:0], 7'h04};
  zdLLziMainzidev5  zdLLziMainzidev5R4 (gzdLLziMainzidev5R4[106:7], gzdLLziMainzidev5R4[6:0], callResR104);
  assign gzdLLziMainzidev5R5 = {gMainzidev[99:0], 7'h05};
  zdLLziMainzidev5  zdLLziMainzidev5R5 (gzdLLziMainzidev5R5[106:7], gzdLLziMainzidev5R5[6:0], callResR105);
  assign gzdLLziMainzidev5R6 = {gMainzidev[99:0], 7'h06};
  zdLLziMainzidev5  zdLLziMainzidev5R6 (gzdLLziMainzidev5R6[106:7], gzdLLziMainzidev5R6[6:0], callResR106);
  assign gzdLLziMainzidev5R7 = {gMainzidev[99:0], 7'h07};
  zdLLziMainzidev5  zdLLziMainzidev5R7 (gzdLLziMainzidev5R7[106:7], gzdLLziMainzidev5R7[6:0], callResR107);
  assign gzdLLziMainzidev5R8 = {gMainzidev[99:0], 7'h08};
  zdLLziMainzidev5  zdLLziMainzidev5R8 (gzdLLziMainzidev5R8[106:7], gzdLLziMainzidev5R8[6:0], callResR108);
  assign gzdLLziMainzidev5R9 = {gMainzidev[99:0], 7'h09};
  zdLLziMainzidev5  zdLLziMainzidev5R9 (gzdLLziMainzidev5R9[106:7], gzdLLziMainzidev5R9[6:0], callResR109);
  assign gzdLLziMainzidev5R10 = {gMainzidev[99:0], 7'h0a};
  zdLLziMainzidev5  zdLLziMainzidev5R10 (gzdLLziMainzidev5R10[106:7], gzdLLziMainzidev5R10[6:0], callResR110);
  assign gzdLLziMainzidev5R11 = {gMainzidev[99:0], 7'h0b};
  zdLLziMainzidev5  zdLLziMainzidev5R11 (gzdLLziMainzidev5R11[106:7], gzdLLziMainzidev5R11[6:0], callResR111);
  assign gzdLLziMainzidev5R12 = {gMainzidev[99:0], 7'h0c};
  zdLLziMainzidev5  zdLLziMainzidev5R12 (gzdLLziMainzidev5R12[106:7], gzdLLziMainzidev5R12[6:0], callResR112);
  assign gzdLLziMainzidev5R13 = {gMainzidev[99:0], 7'h0d};
  zdLLziMainzidev5  zdLLziMainzidev5R13 (gzdLLziMainzidev5R13[106:7], gzdLLziMainzidev5R13[6:0], callResR113);
  assign gzdLLziMainzidev5R14 = {gMainzidev[99:0], 7'h0e};
  zdLLziMainzidev5  zdLLziMainzidev5R14 (gzdLLziMainzidev5R14[106:7], gzdLLziMainzidev5R14[6:0], callResR114);
  assign gzdLLziMainzidev5R15 = {gMainzidev[99:0], 7'h0f};
  zdLLziMainzidev5  zdLLziMainzidev5R15 (gzdLLziMainzidev5R15[106:7], gzdLLziMainzidev5R15[6:0], callResR115);
  assign gzdLLziMainzidev5R16 = {gMainzidev[99:0], 7'h10};
  zdLLziMainzidev5  zdLLziMainzidev5R16 (gzdLLziMainzidev5R16[106:7], gzdLLziMainzidev5R16[6:0], callResR116);
  assign gzdLLziMainzidev5R17 = {gMainzidev[99:0], 7'h11};
  zdLLziMainzidev5  zdLLziMainzidev5R17 (gzdLLziMainzidev5R17[106:7], gzdLLziMainzidev5R17[6:0], callResR117);
  assign gzdLLziMainzidev5R18 = {gMainzidev[99:0], 7'h12};
  zdLLziMainzidev5  zdLLziMainzidev5R18 (gzdLLziMainzidev5R18[106:7], gzdLLziMainzidev5R18[6:0], callResR118);
  assign gzdLLziMainzidev5R19 = {gMainzidev[99:0], 7'h13};
  zdLLziMainzidev5  zdLLziMainzidev5R19 (gzdLLziMainzidev5R19[106:7], gzdLLziMainzidev5R19[6:0], callResR119);
  assign gzdLLziMainzidev5R20 = {gMainzidev[99:0], 7'h14};
  zdLLziMainzidev5  zdLLziMainzidev5R20 (gzdLLziMainzidev5R20[106:7], gzdLLziMainzidev5R20[6:0], callResR120);
  assign gzdLLziMainzidev5R21 = {gMainzidev[99:0], 7'h15};
  zdLLziMainzidev5  zdLLziMainzidev5R21 (gzdLLziMainzidev5R21[106:7], gzdLLziMainzidev5R21[6:0], callResR121);
  assign gzdLLziMainzidev5R22 = {gMainzidev[99:0], 7'h16};
  zdLLziMainzidev5  zdLLziMainzidev5R22 (gzdLLziMainzidev5R22[106:7], gzdLLziMainzidev5R22[6:0], callResR122);
  assign gzdLLziMainzidev5R23 = {gMainzidev[99:0], 7'h17};
  zdLLziMainzidev5  zdLLziMainzidev5R23 (gzdLLziMainzidev5R23[106:7], gzdLLziMainzidev5R23[6:0], callResR123);
  assign gzdLLziMainzidev5R24 = {gMainzidev[99:0], 7'h18};
  zdLLziMainzidev5  zdLLziMainzidev5R24 (gzdLLziMainzidev5R24[106:7], gzdLLziMainzidev5R24[6:0], callResR124);
  assign gzdLLziMainzidev5R25 = {gMainzidev[99:0], 7'h19};
  zdLLziMainzidev5  zdLLziMainzidev5R25 (gzdLLziMainzidev5R25[106:7], gzdLLziMainzidev5R25[6:0], callResR125);
  assign gzdLLziMainzidev5R26 = {gMainzidev[99:0], 7'h1a};
  zdLLziMainzidev5  zdLLziMainzidev5R26 (gzdLLziMainzidev5R26[106:7], gzdLLziMainzidev5R26[6:0], callResR126);
  assign gzdLLziMainzidev5R27 = {gMainzidev[99:0], 7'h1b};
  zdLLziMainzidev5  zdLLziMainzidev5R27 (gzdLLziMainzidev5R27[106:7], gzdLLziMainzidev5R27[6:0], callResR127);
  assign gzdLLziMainzidev5R28 = {gMainzidev[99:0], 7'h1c};
  zdLLziMainzidev5  zdLLziMainzidev5R28 (gzdLLziMainzidev5R28[106:7], gzdLLziMainzidev5R28[6:0], callResR128);
  assign gzdLLziMainzidev5R29 = {gMainzidev[99:0], 7'h1d};
  zdLLziMainzidev5  zdLLziMainzidev5R29 (gzdLLziMainzidev5R29[106:7], gzdLLziMainzidev5R29[6:0], callResR129);
  assign gzdLLziMainzidev5R30 = {gMainzidev[99:0], 7'h1e};
  zdLLziMainzidev5  zdLLziMainzidev5R30 (gzdLLziMainzidev5R30[106:7], gzdLLziMainzidev5R30[6:0], callResR130);
  assign gzdLLziMainzidev5R31 = {gMainzidev[99:0], 7'h1f};
  zdLLziMainzidev5  zdLLziMainzidev5R31 (gzdLLziMainzidev5R31[106:7], gzdLLziMainzidev5R31[6:0], callResR131);
  assign gzdLLziMainzidev5R32 = {gMainzidev[99:0], 7'h20};
  zdLLziMainzidev5  zdLLziMainzidev5R32 (gzdLLziMainzidev5R32[106:7], gzdLLziMainzidev5R32[6:0], callResR132);
  assign gzdLLziMainzidev5R33 = {gMainzidev[99:0], 7'h21};
  zdLLziMainzidev5  zdLLziMainzidev5R33 (gzdLLziMainzidev5R33[106:7], gzdLLziMainzidev5R33[6:0], callResR133);
  assign gzdLLziMainzidev5R34 = {gMainzidev[99:0], 7'h22};
  zdLLziMainzidev5  zdLLziMainzidev5R34 (gzdLLziMainzidev5R34[106:7], gzdLLziMainzidev5R34[6:0], callResR134);
  assign gzdLLziMainzidev5R35 = {gMainzidev[99:0], 7'h23};
  zdLLziMainzidev5  zdLLziMainzidev5R35 (gzdLLziMainzidev5R35[106:7], gzdLLziMainzidev5R35[6:0], callResR135);
  assign gzdLLziMainzidev5R36 = {gMainzidev[99:0], 7'h24};
  zdLLziMainzidev5  zdLLziMainzidev5R36 (gzdLLziMainzidev5R36[106:7], gzdLLziMainzidev5R36[6:0], callResR136);
  assign gzdLLziMainzidev5R37 = {gMainzidev[99:0], 7'h25};
  zdLLziMainzidev5  zdLLziMainzidev5R37 (gzdLLziMainzidev5R37[106:7], gzdLLziMainzidev5R37[6:0], callResR137);
  assign gzdLLziMainzidev5R38 = {gMainzidev[99:0], 7'h26};
  zdLLziMainzidev5  zdLLziMainzidev5R38 (gzdLLziMainzidev5R38[106:7], gzdLLziMainzidev5R38[6:0], callResR138);
  assign gzdLLziMainzidev5R39 = {gMainzidev[99:0], 7'h27};
  zdLLziMainzidev5  zdLLziMainzidev5R39 (gzdLLziMainzidev5R39[106:7], gzdLLziMainzidev5R39[6:0], callResR139);
  assign gzdLLziMainzidev5R40 = {gMainzidev[99:0], 7'h28};
  zdLLziMainzidev5  zdLLziMainzidev5R40 (gzdLLziMainzidev5R40[106:7], gzdLLziMainzidev5R40[6:0], callResR140);
  assign gzdLLziMainzidev5R41 = {gMainzidev[99:0], 7'h29};
  zdLLziMainzidev5  zdLLziMainzidev5R41 (gzdLLziMainzidev5R41[106:7], gzdLLziMainzidev5R41[6:0], callResR141);
  assign gzdLLziMainzidev5R42 = {gMainzidev[99:0], 7'h2a};
  zdLLziMainzidev5  zdLLziMainzidev5R42 (gzdLLziMainzidev5R42[106:7], gzdLLziMainzidev5R42[6:0], callResR142);
  assign gzdLLziMainzidev5R43 = {gMainzidev[99:0], 7'h2b};
  zdLLziMainzidev5  zdLLziMainzidev5R43 (gzdLLziMainzidev5R43[106:7], gzdLLziMainzidev5R43[6:0], callResR143);
  assign gzdLLziMainzidev5R44 = {gMainzidev[99:0], 7'h2c};
  zdLLziMainzidev5  zdLLziMainzidev5R44 (gzdLLziMainzidev5R44[106:7], gzdLLziMainzidev5R44[6:0], callResR144);
  assign gzdLLziMainzidev5R45 = {gMainzidev[99:0], 7'h2d};
  zdLLziMainzidev5  zdLLziMainzidev5R45 (gzdLLziMainzidev5R45[106:7], gzdLLziMainzidev5R45[6:0], callResR145);
  assign gzdLLziMainzidev5R46 = {gMainzidev[99:0], 7'h2e};
  zdLLziMainzidev5  zdLLziMainzidev5R46 (gzdLLziMainzidev5R46[106:7], gzdLLziMainzidev5R46[6:0], callResR146);
  assign gzdLLziMainzidev5R47 = {gMainzidev[99:0], 7'h2f};
  zdLLziMainzidev5  zdLLziMainzidev5R47 (gzdLLziMainzidev5R47[106:7], gzdLLziMainzidev5R47[6:0], callResR147);
  assign gzdLLziMainzidev5R48 = {gMainzidev[99:0], 7'h30};
  zdLLziMainzidev5  zdLLziMainzidev5R48 (gzdLLziMainzidev5R48[106:7], gzdLLziMainzidev5R48[6:0], callResR148);
  assign gzdLLziMainzidev5R49 = {gMainzidev[99:0], 7'h31};
  zdLLziMainzidev5  zdLLziMainzidev5R49 (gzdLLziMainzidev5R49[106:7], gzdLLziMainzidev5R49[6:0], callResR149);
  assign gzdLLziMainzidev5R50 = {gMainzidev[99:0], 7'h32};
  zdLLziMainzidev5  zdLLziMainzidev5R50 (gzdLLziMainzidev5R50[106:7], gzdLLziMainzidev5R50[6:0], callResR150);
  assign gzdLLziMainzidev5R51 = {gMainzidev[99:0], 7'h33};
  zdLLziMainzidev5  zdLLziMainzidev5R51 (gzdLLziMainzidev5R51[106:7], gzdLLziMainzidev5R51[6:0], callResR151);
  assign gzdLLziMainzidev5R52 = {gMainzidev[99:0], 7'h34};
  zdLLziMainzidev5  zdLLziMainzidev5R52 (gzdLLziMainzidev5R52[106:7], gzdLLziMainzidev5R52[6:0], callResR152);
  assign gzdLLziMainzidev5R53 = {gMainzidev[99:0], 7'h35};
  zdLLziMainzidev5  zdLLziMainzidev5R53 (gzdLLziMainzidev5R53[106:7], gzdLLziMainzidev5R53[6:0], callResR153);
  assign gzdLLziMainzidev5R54 = {gMainzidev[99:0], 7'h36};
  zdLLziMainzidev5  zdLLziMainzidev5R54 (gzdLLziMainzidev5R54[106:7], gzdLLziMainzidev5R54[6:0], callResR154);
  assign gzdLLziMainzidev5R55 = {gMainzidev[99:0], 7'h37};
  zdLLziMainzidev5  zdLLziMainzidev5R55 (gzdLLziMainzidev5R55[106:7], gzdLLziMainzidev5R55[6:0], callResR155);
  assign gzdLLziMainzidev5R56 = {gMainzidev[99:0], 7'h38};
  zdLLziMainzidev5  zdLLziMainzidev5R56 (gzdLLziMainzidev5R56[106:7], gzdLLziMainzidev5R56[6:0], callResR156);
  assign gzdLLziMainzidev5R57 = {gMainzidev[99:0], 7'h39};
  zdLLziMainzidev5  zdLLziMainzidev5R57 (gzdLLziMainzidev5R57[106:7], gzdLLziMainzidev5R57[6:0], callResR157);
  assign gzdLLziMainzidev5R58 = {gMainzidev[99:0], 7'h3a};
  zdLLziMainzidev5  zdLLziMainzidev5R58 (gzdLLziMainzidev5R58[106:7], gzdLLziMainzidev5R58[6:0], callResR158);
  assign gzdLLziMainzidev5R59 = {gMainzidev[99:0], 7'h3b};
  zdLLziMainzidev5  zdLLziMainzidev5R59 (gzdLLziMainzidev5R59[106:7], gzdLLziMainzidev5R59[6:0], callResR159);
  assign gzdLLziMainzidev5R60 = {gMainzidev[99:0], 7'h3c};
  zdLLziMainzidev5  zdLLziMainzidev5R60 (gzdLLziMainzidev5R60[106:7], gzdLLziMainzidev5R60[6:0], callResR160);
  assign gzdLLziMainzidev5R61 = {gMainzidev[99:0], 7'h3d};
  zdLLziMainzidev5  zdLLziMainzidev5R61 (gzdLLziMainzidev5R61[106:7], gzdLLziMainzidev5R61[6:0], callResR161);
  assign gzdLLziMainzidev5R62 = {gMainzidev[99:0], 7'h3e};
  zdLLziMainzidev5  zdLLziMainzidev5R62 (gzdLLziMainzidev5R62[106:7], gzdLLziMainzidev5R62[6:0], callResR162);
  assign gzdLLziMainzidev5R63 = {gMainzidev[99:0], 7'h3f};
  zdLLziMainzidev5  zdLLziMainzidev5R63 (gzdLLziMainzidev5R63[106:7], gzdLLziMainzidev5R63[6:0], callResR163);
  assign gzdLLziMainzidev5R64 = {gMainzidev[99:0], 7'h40};
  zdLLziMainzidev5  zdLLziMainzidev5R64 (gzdLLziMainzidev5R64[106:7], gzdLLziMainzidev5R64[6:0], callResR164);
  assign gzdLLziMainzidev5R65 = {gMainzidev[99:0], 7'h41};
  zdLLziMainzidev5  zdLLziMainzidev5R65 (gzdLLziMainzidev5R65[106:7], gzdLLziMainzidev5R65[6:0], callResR165);
  assign gzdLLziMainzidev5R66 = {gMainzidev[99:0], 7'h42};
  zdLLziMainzidev5  zdLLziMainzidev5R66 (gzdLLziMainzidev5R66[106:7], gzdLLziMainzidev5R66[6:0], callResR166);
  assign gzdLLziMainzidev5R67 = {gMainzidev[99:0], 7'h43};
  zdLLziMainzidev5  zdLLziMainzidev5R67 (gzdLLziMainzidev5R67[106:7], gzdLLziMainzidev5R67[6:0], callResR167);
  assign gzdLLziMainzidev5R68 = {gMainzidev[99:0], 7'h44};
  zdLLziMainzidev5  zdLLziMainzidev5R68 (gzdLLziMainzidev5R68[106:7], gzdLLziMainzidev5R68[6:0], callResR168);
  assign gzdLLziMainzidev5R69 = {gMainzidev[99:0], 7'h45};
  zdLLziMainzidev5  zdLLziMainzidev5R69 (gzdLLziMainzidev5R69[106:7], gzdLLziMainzidev5R69[6:0], callResR169);
  assign gzdLLziMainzidev5R70 = {gMainzidev[99:0], 7'h46};
  zdLLziMainzidev5  zdLLziMainzidev5R70 (gzdLLziMainzidev5R70[106:7], gzdLLziMainzidev5R70[6:0], callResR170);
  assign gzdLLziMainzidev5R71 = {gMainzidev[99:0], 7'h47};
  zdLLziMainzidev5  zdLLziMainzidev5R71 (gzdLLziMainzidev5R71[106:7], gzdLLziMainzidev5R71[6:0], callResR171);
  assign gzdLLziMainzidev5R72 = {gMainzidev[99:0], 7'h48};
  zdLLziMainzidev5  zdLLziMainzidev5R72 (gzdLLziMainzidev5R72[106:7], gzdLLziMainzidev5R72[6:0], callResR172);
  assign gzdLLziMainzidev5R73 = {gMainzidev[99:0], 7'h49};
  zdLLziMainzidev5  zdLLziMainzidev5R73 (gzdLLziMainzidev5R73[106:7], gzdLLziMainzidev5R73[6:0], callResR173);
  assign gzdLLziMainzidev5R74 = {gMainzidev[99:0], 7'h4a};
  zdLLziMainzidev5  zdLLziMainzidev5R74 (gzdLLziMainzidev5R74[106:7], gzdLLziMainzidev5R74[6:0], callResR174);
  assign gzdLLziMainzidev5R75 = {gMainzidev[99:0], 7'h4b};
  zdLLziMainzidev5  zdLLziMainzidev5R75 (gzdLLziMainzidev5R75[106:7], gzdLLziMainzidev5R75[6:0], callResR175);
  assign gzdLLziMainzidev5R76 = {gMainzidev[99:0], 7'h4c};
  zdLLziMainzidev5  zdLLziMainzidev5R76 (gzdLLziMainzidev5R76[106:7], gzdLLziMainzidev5R76[6:0], callResR176);
  assign gzdLLziMainzidev5R77 = {gMainzidev[99:0], 7'h4d};
  zdLLziMainzidev5  zdLLziMainzidev5R77 (gzdLLziMainzidev5R77[106:7], gzdLLziMainzidev5R77[6:0], callResR177);
  assign gzdLLziMainzidev5R78 = {gMainzidev[99:0], 7'h4e};
  zdLLziMainzidev5  zdLLziMainzidev5R78 (gzdLLziMainzidev5R78[106:7], gzdLLziMainzidev5R78[6:0], callResR178);
  assign gzdLLziMainzidev5R79 = {gMainzidev[99:0], 7'h4f};
  zdLLziMainzidev5  zdLLziMainzidev5R79 (gzdLLziMainzidev5R79[106:7], gzdLLziMainzidev5R79[6:0], callResR179);
  assign gzdLLziMainzidev5R80 = {gMainzidev[99:0], 7'h50};
  zdLLziMainzidev5  zdLLziMainzidev5R80 (gzdLLziMainzidev5R80[106:7], gzdLLziMainzidev5R80[6:0], callResR180);
  assign gzdLLziMainzidev5R81 = {gMainzidev[99:0], 7'h51};
  zdLLziMainzidev5  zdLLziMainzidev5R81 (gzdLLziMainzidev5R81[106:7], gzdLLziMainzidev5R81[6:0], callResR181);
  assign gzdLLziMainzidev5R82 = {gMainzidev[99:0], 7'h52};
  zdLLziMainzidev5  zdLLziMainzidev5R82 (gzdLLziMainzidev5R82[106:7], gzdLLziMainzidev5R82[6:0], callResR182);
  assign gzdLLziMainzidev5R83 = {gMainzidev[99:0], 7'h53};
  zdLLziMainzidev5  zdLLziMainzidev5R83 (gzdLLziMainzidev5R83[106:7], gzdLLziMainzidev5R83[6:0], callResR183);
  assign gzdLLziMainzidev5R84 = {gMainzidev[99:0], 7'h54};
  zdLLziMainzidev5  zdLLziMainzidev5R84 (gzdLLziMainzidev5R84[106:7], gzdLLziMainzidev5R84[6:0], callResR184);
  assign gzdLLziMainzidev5R85 = {gMainzidev[99:0], 7'h55};
  zdLLziMainzidev5  zdLLziMainzidev5R85 (gzdLLziMainzidev5R85[106:7], gzdLLziMainzidev5R85[6:0], callResR185);
  assign gzdLLziMainzidev5R86 = {gMainzidev[99:0], 7'h56};
  zdLLziMainzidev5  zdLLziMainzidev5R86 (gzdLLziMainzidev5R86[106:7], gzdLLziMainzidev5R86[6:0], callResR186);
  assign gzdLLziMainzidev5R87 = {gMainzidev[99:0], 7'h57};
  zdLLziMainzidev5  zdLLziMainzidev5R87 (gzdLLziMainzidev5R87[106:7], gzdLLziMainzidev5R87[6:0], callResR187);
  assign gzdLLziMainzidev5R88 = {gMainzidev[99:0], 7'h58};
  zdLLziMainzidev5  zdLLziMainzidev5R88 (gzdLLziMainzidev5R88[106:7], gzdLLziMainzidev5R88[6:0], callResR188);
  assign gzdLLziMainzidev5R89 = {gMainzidev[99:0], 7'h59};
  zdLLziMainzidev5  zdLLziMainzidev5R89 (gzdLLziMainzidev5R89[106:7], gzdLLziMainzidev5R89[6:0], callResR189);
  assign gzdLLziMainzidev5R90 = {gMainzidev[99:0], 7'h5a};
  zdLLziMainzidev5  zdLLziMainzidev5R90 (gzdLLziMainzidev5R90[106:7], gzdLLziMainzidev5R90[6:0], callResR190);
  assign gzdLLziMainzidev5R91 = {gMainzidev[99:0], 7'h5b};
  zdLLziMainzidev5  zdLLziMainzidev5R91 (gzdLLziMainzidev5R91[106:7], gzdLLziMainzidev5R91[6:0], callResR191);
  assign gzdLLziMainzidev5R92 = {gMainzidev[99:0], 7'h5c};
  zdLLziMainzidev5  zdLLziMainzidev5R92 (gzdLLziMainzidev5R92[106:7], gzdLLziMainzidev5R92[6:0], callResR192);
  assign gzdLLziMainzidev5R93 = {gMainzidev[99:0], 7'h5d};
  zdLLziMainzidev5  zdLLziMainzidev5R93 (gzdLLziMainzidev5R93[106:7], gzdLLziMainzidev5R93[6:0], callResR193);
  assign gzdLLziMainzidev5R94 = {gMainzidev[99:0], 7'h5e};
  zdLLziMainzidev5  zdLLziMainzidev5R94 (gzdLLziMainzidev5R94[106:7], gzdLLziMainzidev5R94[6:0], callResR194);
  assign gzdLLziMainzidev5R95 = {gMainzidev[99:0], 7'h5f};
  zdLLziMainzidev5  zdLLziMainzidev5R95 (gzdLLziMainzidev5R95[106:7], gzdLLziMainzidev5R95[6:0], callResR195);
  assign gzdLLziMainzidev5R96 = {gMainzidev[99:0], 7'h60};
  zdLLziMainzidev5  zdLLziMainzidev5R96 (gzdLLziMainzidev5R96[106:7], gzdLLziMainzidev5R96[6:0], callResR196);
  assign gzdLLziMainzidev5R97 = {gMainzidev[99:0], 7'h61};
  zdLLziMainzidev5  zdLLziMainzidev5R97 (gzdLLziMainzidev5R97[106:7], gzdLLziMainzidev5R97[6:0], callResR197);
  assign gzdLLziMainzidev5R98 = {gMainzidev[99:0], 7'h62};
  zdLLziMainzidev5  zdLLziMainzidev5R98 (gzdLLziMainzidev5R98[106:7], gzdLLziMainzidev5R98[6:0], callResR198);
  assign gzdLLziMainzidev5R99 = {gMainzidev[99:0], 7'h63};
  zdLLziMainzidev5  zdLLziMainzidev5R99 (gzdLLziMainzidev5R99[106:7], gzdLLziMainzidev5R99[6:0], callResR199);
  assign gzdLLziMainzidev8 = {gMainzidev[99:0], 7'h00};
  zdLLziMainzidev8  zdLLziMainzidev8 (gzdLLziMainzidev8[106:7], gzdLLziMainzidev8[6:0], callResR200);
  assign gzdLLziMainzidev8R1 = {gMainzidev[99:0], 7'h01};
  zdLLziMainzidev8  zdLLziMainzidev8R1 (gzdLLziMainzidev8R1[106:7], gzdLLziMainzidev8R1[6:0], callResR201);
  assign gzdLLziMainzidev8R2 = {gMainzidev[99:0], 7'h02};
  zdLLziMainzidev8  zdLLziMainzidev8R2 (gzdLLziMainzidev8R2[106:7], gzdLLziMainzidev8R2[6:0], callResR202);
  assign gzdLLziMainzidev8R3 = {gMainzidev[99:0], 7'h03};
  zdLLziMainzidev8  zdLLziMainzidev8R3 (gzdLLziMainzidev8R3[106:7], gzdLLziMainzidev8R3[6:0], callResR203);
  assign gzdLLziMainzidev8R4 = {gMainzidev[99:0], 7'h04};
  zdLLziMainzidev8  zdLLziMainzidev8R4 (gzdLLziMainzidev8R4[106:7], gzdLLziMainzidev8R4[6:0], callResR204);
  assign gzdLLziMainzidev8R5 = {gMainzidev[99:0], 7'h05};
  zdLLziMainzidev8  zdLLziMainzidev8R5 (gzdLLziMainzidev8R5[106:7], gzdLLziMainzidev8R5[6:0], callResR205);
  assign gzdLLziMainzidev8R6 = {gMainzidev[99:0], 7'h06};
  zdLLziMainzidev8  zdLLziMainzidev8R6 (gzdLLziMainzidev8R6[106:7], gzdLLziMainzidev8R6[6:0], callResR206);
  assign gzdLLziMainzidev8R7 = {gMainzidev[99:0], 7'h07};
  zdLLziMainzidev8  zdLLziMainzidev8R7 (gzdLLziMainzidev8R7[106:7], gzdLLziMainzidev8R7[6:0], callResR207);
  assign gzdLLziMainzidev8R8 = {gMainzidev[99:0], 7'h08};
  zdLLziMainzidev8  zdLLziMainzidev8R8 (gzdLLziMainzidev8R8[106:7], gzdLLziMainzidev8R8[6:0], callResR208);
  assign gzdLLziMainzidev8R9 = {gMainzidev[99:0], 7'h09};
  zdLLziMainzidev8  zdLLziMainzidev8R9 (gzdLLziMainzidev8R9[106:7], gzdLLziMainzidev8R9[6:0], callResR209);
  assign gzdLLziMainzidev8R10 = {gMainzidev[99:0], 7'h0a};
  zdLLziMainzidev8  zdLLziMainzidev8R10 (gzdLLziMainzidev8R10[106:7], gzdLLziMainzidev8R10[6:0], callResR210);
  assign gzdLLziMainzidev8R11 = {gMainzidev[99:0], 7'h0b};
  zdLLziMainzidev8  zdLLziMainzidev8R11 (gzdLLziMainzidev8R11[106:7], gzdLLziMainzidev8R11[6:0], callResR211);
  assign gzdLLziMainzidev8R12 = {gMainzidev[99:0], 7'h0c};
  zdLLziMainzidev8  zdLLziMainzidev8R12 (gzdLLziMainzidev8R12[106:7], gzdLLziMainzidev8R12[6:0], callResR212);
  assign gzdLLziMainzidev8R13 = {gMainzidev[99:0], 7'h0d};
  zdLLziMainzidev8  zdLLziMainzidev8R13 (gzdLLziMainzidev8R13[106:7], gzdLLziMainzidev8R13[6:0], callResR213);
  assign gzdLLziMainzidev8R14 = {gMainzidev[99:0], 7'h0e};
  zdLLziMainzidev8  zdLLziMainzidev8R14 (gzdLLziMainzidev8R14[106:7], gzdLLziMainzidev8R14[6:0], callResR214);
  assign gzdLLziMainzidev8R15 = {gMainzidev[99:0], 7'h0f};
  zdLLziMainzidev8  zdLLziMainzidev8R15 (gzdLLziMainzidev8R15[106:7], gzdLLziMainzidev8R15[6:0], callResR215);
  assign gzdLLziMainzidev8R16 = {gMainzidev[99:0], 7'h10};
  zdLLziMainzidev8  zdLLziMainzidev8R16 (gzdLLziMainzidev8R16[106:7], gzdLLziMainzidev8R16[6:0], callResR216);
  assign gzdLLziMainzidev8R17 = {gMainzidev[99:0], 7'h11};
  zdLLziMainzidev8  zdLLziMainzidev8R17 (gzdLLziMainzidev8R17[106:7], gzdLLziMainzidev8R17[6:0], callResR217);
  assign gzdLLziMainzidev8R18 = {gMainzidev[99:0], 7'h12};
  zdLLziMainzidev8  zdLLziMainzidev8R18 (gzdLLziMainzidev8R18[106:7], gzdLLziMainzidev8R18[6:0], callResR218);
  assign gzdLLziMainzidev8R19 = {gMainzidev[99:0], 7'h13};
  zdLLziMainzidev8  zdLLziMainzidev8R19 (gzdLLziMainzidev8R19[106:7], gzdLLziMainzidev8R19[6:0], callResR219);
  assign gzdLLziMainzidev8R20 = {gMainzidev[99:0], 7'h14};
  zdLLziMainzidev8  zdLLziMainzidev8R20 (gzdLLziMainzidev8R20[106:7], gzdLLziMainzidev8R20[6:0], callResR220);
  assign gzdLLziMainzidev8R21 = {gMainzidev[99:0], 7'h15};
  zdLLziMainzidev8  zdLLziMainzidev8R21 (gzdLLziMainzidev8R21[106:7], gzdLLziMainzidev8R21[6:0], callResR221);
  assign gzdLLziMainzidev8R22 = {gMainzidev[99:0], 7'h16};
  zdLLziMainzidev8  zdLLziMainzidev8R22 (gzdLLziMainzidev8R22[106:7], gzdLLziMainzidev8R22[6:0], callResR222);
  assign gzdLLziMainzidev8R23 = {gMainzidev[99:0], 7'h17};
  zdLLziMainzidev8  zdLLziMainzidev8R23 (gzdLLziMainzidev8R23[106:7], gzdLLziMainzidev8R23[6:0], callResR223);
  assign gzdLLziMainzidev8R24 = {gMainzidev[99:0], 7'h18};
  zdLLziMainzidev8  zdLLziMainzidev8R24 (gzdLLziMainzidev8R24[106:7], gzdLLziMainzidev8R24[6:0], callResR224);
  assign gzdLLziMainzidev8R25 = {gMainzidev[99:0], 7'h19};
  zdLLziMainzidev8  zdLLziMainzidev8R25 (gzdLLziMainzidev8R25[106:7], gzdLLziMainzidev8R25[6:0], callResR225);
  assign gzdLLziMainzidev8R26 = {gMainzidev[99:0], 7'h1a};
  zdLLziMainzidev8  zdLLziMainzidev8R26 (gzdLLziMainzidev8R26[106:7], gzdLLziMainzidev8R26[6:0], callResR226);
  assign gzdLLziMainzidev8R27 = {gMainzidev[99:0], 7'h1b};
  zdLLziMainzidev8  zdLLziMainzidev8R27 (gzdLLziMainzidev8R27[106:7], gzdLLziMainzidev8R27[6:0], callResR227);
  assign gzdLLziMainzidev8R28 = {gMainzidev[99:0], 7'h1c};
  zdLLziMainzidev8  zdLLziMainzidev8R28 (gzdLLziMainzidev8R28[106:7], gzdLLziMainzidev8R28[6:0], callResR228);
  assign gzdLLziMainzidev8R29 = {gMainzidev[99:0], 7'h1d};
  zdLLziMainzidev8  zdLLziMainzidev8R29 (gzdLLziMainzidev8R29[106:7], gzdLLziMainzidev8R29[6:0], callResR229);
  assign gzdLLziMainzidev8R30 = {gMainzidev[99:0], 7'h1e};
  zdLLziMainzidev8  zdLLziMainzidev8R30 (gzdLLziMainzidev8R30[106:7], gzdLLziMainzidev8R30[6:0], callResR230);
  assign gzdLLziMainzidev8R31 = {gMainzidev[99:0], 7'h1f};
  zdLLziMainzidev8  zdLLziMainzidev8R31 (gzdLLziMainzidev8R31[106:7], gzdLLziMainzidev8R31[6:0], callResR231);
  assign gzdLLziMainzidev8R32 = {gMainzidev[99:0], 7'h20};
  zdLLziMainzidev8  zdLLziMainzidev8R32 (gzdLLziMainzidev8R32[106:7], gzdLLziMainzidev8R32[6:0], callResR232);
  assign gzdLLziMainzidev8R33 = {gMainzidev[99:0], 7'h21};
  zdLLziMainzidev8  zdLLziMainzidev8R33 (gzdLLziMainzidev8R33[106:7], gzdLLziMainzidev8R33[6:0], callResR233);
  assign gzdLLziMainzidev8R34 = {gMainzidev[99:0], 7'h22};
  zdLLziMainzidev8  zdLLziMainzidev8R34 (gzdLLziMainzidev8R34[106:7], gzdLLziMainzidev8R34[6:0], callResR234);
  assign gzdLLziMainzidev8R35 = {gMainzidev[99:0], 7'h23};
  zdLLziMainzidev8  zdLLziMainzidev8R35 (gzdLLziMainzidev8R35[106:7], gzdLLziMainzidev8R35[6:0], callResR235);
  assign gzdLLziMainzidev8R36 = {gMainzidev[99:0], 7'h24};
  zdLLziMainzidev8  zdLLziMainzidev8R36 (gzdLLziMainzidev8R36[106:7], gzdLLziMainzidev8R36[6:0], callResR236);
  assign gzdLLziMainzidev8R37 = {gMainzidev[99:0], 7'h25};
  zdLLziMainzidev8  zdLLziMainzidev8R37 (gzdLLziMainzidev8R37[106:7], gzdLLziMainzidev8R37[6:0], callResR237);
  assign gzdLLziMainzidev8R38 = {gMainzidev[99:0], 7'h26};
  zdLLziMainzidev8  zdLLziMainzidev8R38 (gzdLLziMainzidev8R38[106:7], gzdLLziMainzidev8R38[6:0], callResR238);
  assign gzdLLziMainzidev8R39 = {gMainzidev[99:0], 7'h27};
  zdLLziMainzidev8  zdLLziMainzidev8R39 (gzdLLziMainzidev8R39[106:7], gzdLLziMainzidev8R39[6:0], callResR239);
  assign gzdLLziMainzidev8R40 = {gMainzidev[99:0], 7'h28};
  zdLLziMainzidev8  zdLLziMainzidev8R40 (gzdLLziMainzidev8R40[106:7], gzdLLziMainzidev8R40[6:0], callResR240);
  assign gzdLLziMainzidev8R41 = {gMainzidev[99:0], 7'h29};
  zdLLziMainzidev8  zdLLziMainzidev8R41 (gzdLLziMainzidev8R41[106:7], gzdLLziMainzidev8R41[6:0], callResR241);
  assign gzdLLziMainzidev8R42 = {gMainzidev[99:0], 7'h2a};
  zdLLziMainzidev8  zdLLziMainzidev8R42 (gzdLLziMainzidev8R42[106:7], gzdLLziMainzidev8R42[6:0], callResR242);
  assign gzdLLziMainzidev8R43 = {gMainzidev[99:0], 7'h2b};
  zdLLziMainzidev8  zdLLziMainzidev8R43 (gzdLLziMainzidev8R43[106:7], gzdLLziMainzidev8R43[6:0], callResR243);
  assign gzdLLziMainzidev8R44 = {gMainzidev[99:0], 7'h2c};
  zdLLziMainzidev8  zdLLziMainzidev8R44 (gzdLLziMainzidev8R44[106:7], gzdLLziMainzidev8R44[6:0], callResR244);
  assign gzdLLziMainzidev8R45 = {gMainzidev[99:0], 7'h2d};
  zdLLziMainzidev8  zdLLziMainzidev8R45 (gzdLLziMainzidev8R45[106:7], gzdLLziMainzidev8R45[6:0], callResR245);
  assign gzdLLziMainzidev8R46 = {gMainzidev[99:0], 7'h2e};
  zdLLziMainzidev8  zdLLziMainzidev8R46 (gzdLLziMainzidev8R46[106:7], gzdLLziMainzidev8R46[6:0], callResR246);
  assign gzdLLziMainzidev8R47 = {gMainzidev[99:0], 7'h2f};
  zdLLziMainzidev8  zdLLziMainzidev8R47 (gzdLLziMainzidev8R47[106:7], gzdLLziMainzidev8R47[6:0], callResR247);
  assign gzdLLziMainzidev8R48 = {gMainzidev[99:0], 7'h30};
  zdLLziMainzidev8  zdLLziMainzidev8R48 (gzdLLziMainzidev8R48[106:7], gzdLLziMainzidev8R48[6:0], callResR248);
  assign gzdLLziMainzidev8R49 = {gMainzidev[99:0], 7'h31};
  zdLLziMainzidev8  zdLLziMainzidev8R49 (gzdLLziMainzidev8R49[106:7], gzdLLziMainzidev8R49[6:0], callResR249);
  assign gzdLLziMainzidev8R50 = {gMainzidev[99:0], 7'h32};
  zdLLziMainzidev8  zdLLziMainzidev8R50 (gzdLLziMainzidev8R50[106:7], gzdLLziMainzidev8R50[6:0], callResR250);
  assign gzdLLziMainzidev8R51 = {gMainzidev[99:0], 7'h33};
  zdLLziMainzidev8  zdLLziMainzidev8R51 (gzdLLziMainzidev8R51[106:7], gzdLLziMainzidev8R51[6:0], callResR251);
  assign gzdLLziMainzidev8R52 = {gMainzidev[99:0], 7'h34};
  zdLLziMainzidev8  zdLLziMainzidev8R52 (gzdLLziMainzidev8R52[106:7], gzdLLziMainzidev8R52[6:0], callResR252);
  assign gzdLLziMainzidev8R53 = {gMainzidev[99:0], 7'h35};
  zdLLziMainzidev8  zdLLziMainzidev8R53 (gzdLLziMainzidev8R53[106:7], gzdLLziMainzidev8R53[6:0], callResR253);
  assign gzdLLziMainzidev8R54 = {gMainzidev[99:0], 7'h36};
  zdLLziMainzidev8  zdLLziMainzidev8R54 (gzdLLziMainzidev8R54[106:7], gzdLLziMainzidev8R54[6:0], callResR254);
  assign gzdLLziMainzidev8R55 = {gMainzidev[99:0], 7'h37};
  zdLLziMainzidev8  zdLLziMainzidev8R55 (gzdLLziMainzidev8R55[106:7], gzdLLziMainzidev8R55[6:0], callResR255);
  assign gzdLLziMainzidev8R56 = {gMainzidev[99:0], 7'h38};
  zdLLziMainzidev8  zdLLziMainzidev8R56 (gzdLLziMainzidev8R56[106:7], gzdLLziMainzidev8R56[6:0], callResR256);
  assign gzdLLziMainzidev8R57 = {gMainzidev[99:0], 7'h39};
  zdLLziMainzidev8  zdLLziMainzidev8R57 (gzdLLziMainzidev8R57[106:7], gzdLLziMainzidev8R57[6:0], callResR257);
  assign gzdLLziMainzidev8R58 = {gMainzidev[99:0], 7'h3a};
  zdLLziMainzidev8  zdLLziMainzidev8R58 (gzdLLziMainzidev8R58[106:7], gzdLLziMainzidev8R58[6:0], callResR258);
  assign gzdLLziMainzidev8R59 = {gMainzidev[99:0], 7'h3b};
  zdLLziMainzidev8  zdLLziMainzidev8R59 (gzdLLziMainzidev8R59[106:7], gzdLLziMainzidev8R59[6:0], callResR259);
  assign gzdLLziMainzidev8R60 = {gMainzidev[99:0], 7'h3c};
  zdLLziMainzidev8  zdLLziMainzidev8R60 (gzdLLziMainzidev8R60[106:7], gzdLLziMainzidev8R60[6:0], callResR260);
  assign gzdLLziMainzidev8R61 = {gMainzidev[99:0], 7'h3d};
  zdLLziMainzidev8  zdLLziMainzidev8R61 (gzdLLziMainzidev8R61[106:7], gzdLLziMainzidev8R61[6:0], callResR261);
  assign gzdLLziMainzidev8R62 = {gMainzidev[99:0], 7'h3e};
  zdLLziMainzidev8  zdLLziMainzidev8R62 (gzdLLziMainzidev8R62[106:7], gzdLLziMainzidev8R62[6:0], callResR262);
  assign gzdLLziMainzidev8R63 = {gMainzidev[99:0], 7'h3f};
  zdLLziMainzidev8  zdLLziMainzidev8R63 (gzdLLziMainzidev8R63[106:7], gzdLLziMainzidev8R63[6:0], callResR263);
  assign gzdLLziMainzidev8R64 = {gMainzidev[99:0], 7'h40};
  zdLLziMainzidev8  zdLLziMainzidev8R64 (gzdLLziMainzidev8R64[106:7], gzdLLziMainzidev8R64[6:0], callResR264);
  assign gzdLLziMainzidev8R65 = {gMainzidev[99:0], 7'h41};
  zdLLziMainzidev8  zdLLziMainzidev8R65 (gzdLLziMainzidev8R65[106:7], gzdLLziMainzidev8R65[6:0], callResR265);
  assign gzdLLziMainzidev8R66 = {gMainzidev[99:0], 7'h42};
  zdLLziMainzidev8  zdLLziMainzidev8R66 (gzdLLziMainzidev8R66[106:7], gzdLLziMainzidev8R66[6:0], callResR266);
  assign gzdLLziMainzidev8R67 = {gMainzidev[99:0], 7'h43};
  zdLLziMainzidev8  zdLLziMainzidev8R67 (gzdLLziMainzidev8R67[106:7], gzdLLziMainzidev8R67[6:0], callResR267);
  assign gzdLLziMainzidev8R68 = {gMainzidev[99:0], 7'h44};
  zdLLziMainzidev8  zdLLziMainzidev8R68 (gzdLLziMainzidev8R68[106:7], gzdLLziMainzidev8R68[6:0], callResR268);
  assign gzdLLziMainzidev8R69 = {gMainzidev[99:0], 7'h45};
  zdLLziMainzidev8  zdLLziMainzidev8R69 (gzdLLziMainzidev8R69[106:7], gzdLLziMainzidev8R69[6:0], callResR269);
  assign gzdLLziMainzidev8R70 = {gMainzidev[99:0], 7'h46};
  zdLLziMainzidev8  zdLLziMainzidev8R70 (gzdLLziMainzidev8R70[106:7], gzdLLziMainzidev8R70[6:0], callResR270);
  assign gzdLLziMainzidev8R71 = {gMainzidev[99:0], 7'h47};
  zdLLziMainzidev8  zdLLziMainzidev8R71 (gzdLLziMainzidev8R71[106:7], gzdLLziMainzidev8R71[6:0], callResR271);
  assign gzdLLziMainzidev8R72 = {gMainzidev[99:0], 7'h48};
  zdLLziMainzidev8  zdLLziMainzidev8R72 (gzdLLziMainzidev8R72[106:7], gzdLLziMainzidev8R72[6:0], callResR272);
  assign gzdLLziMainzidev8R73 = {gMainzidev[99:0], 7'h49};
  zdLLziMainzidev8  zdLLziMainzidev8R73 (gzdLLziMainzidev8R73[106:7], gzdLLziMainzidev8R73[6:0], callResR273);
  assign gzdLLziMainzidev8R74 = {gMainzidev[99:0], 7'h4a};
  zdLLziMainzidev8  zdLLziMainzidev8R74 (gzdLLziMainzidev8R74[106:7], gzdLLziMainzidev8R74[6:0], callResR274);
  assign gzdLLziMainzidev8R75 = {gMainzidev[99:0], 7'h4b};
  zdLLziMainzidev8  zdLLziMainzidev8R75 (gzdLLziMainzidev8R75[106:7], gzdLLziMainzidev8R75[6:0], callResR275);
  assign gzdLLziMainzidev8R76 = {gMainzidev[99:0], 7'h4c};
  zdLLziMainzidev8  zdLLziMainzidev8R76 (gzdLLziMainzidev8R76[106:7], gzdLLziMainzidev8R76[6:0], callResR276);
  assign gzdLLziMainzidev8R77 = {gMainzidev[99:0], 7'h4d};
  zdLLziMainzidev8  zdLLziMainzidev8R77 (gzdLLziMainzidev8R77[106:7], gzdLLziMainzidev8R77[6:0], callResR277);
  assign gzdLLziMainzidev8R78 = {gMainzidev[99:0], 7'h4e};
  zdLLziMainzidev8  zdLLziMainzidev8R78 (gzdLLziMainzidev8R78[106:7], gzdLLziMainzidev8R78[6:0], callResR278);
  assign gzdLLziMainzidev8R79 = {gMainzidev[99:0], 7'h4f};
  zdLLziMainzidev8  zdLLziMainzidev8R79 (gzdLLziMainzidev8R79[106:7], gzdLLziMainzidev8R79[6:0], callResR279);
  assign gzdLLziMainzidev8R80 = {gMainzidev[99:0], 7'h50};
  zdLLziMainzidev8  zdLLziMainzidev8R80 (gzdLLziMainzidev8R80[106:7], gzdLLziMainzidev8R80[6:0], callResR280);
  assign gzdLLziMainzidev8R81 = {gMainzidev[99:0], 7'h51};
  zdLLziMainzidev8  zdLLziMainzidev8R81 (gzdLLziMainzidev8R81[106:7], gzdLLziMainzidev8R81[6:0], callResR281);
  assign gzdLLziMainzidev8R82 = {gMainzidev[99:0], 7'h52};
  zdLLziMainzidev8  zdLLziMainzidev8R82 (gzdLLziMainzidev8R82[106:7], gzdLLziMainzidev8R82[6:0], callResR282);
  assign gzdLLziMainzidev8R83 = {gMainzidev[99:0], 7'h53};
  zdLLziMainzidev8  zdLLziMainzidev8R83 (gzdLLziMainzidev8R83[106:7], gzdLLziMainzidev8R83[6:0], callResR283);
  assign gzdLLziMainzidev8R84 = {gMainzidev[99:0], 7'h54};
  zdLLziMainzidev8  zdLLziMainzidev8R84 (gzdLLziMainzidev8R84[106:7], gzdLLziMainzidev8R84[6:0], callResR284);
  assign gzdLLziMainzidev8R85 = {gMainzidev[99:0], 7'h55};
  zdLLziMainzidev8  zdLLziMainzidev8R85 (gzdLLziMainzidev8R85[106:7], gzdLLziMainzidev8R85[6:0], callResR285);
  assign gzdLLziMainzidev8R86 = {gMainzidev[99:0], 7'h56};
  zdLLziMainzidev8  zdLLziMainzidev8R86 (gzdLLziMainzidev8R86[106:7], gzdLLziMainzidev8R86[6:0], callResR286);
  assign gzdLLziMainzidev8R87 = {gMainzidev[99:0], 7'h57};
  zdLLziMainzidev8  zdLLziMainzidev8R87 (gzdLLziMainzidev8R87[106:7], gzdLLziMainzidev8R87[6:0], callResR287);
  assign gzdLLziMainzidev8R88 = {gMainzidev[99:0], 7'h58};
  zdLLziMainzidev8  zdLLziMainzidev8R88 (gzdLLziMainzidev8R88[106:7], gzdLLziMainzidev8R88[6:0], callResR288);
  assign gzdLLziMainzidev8R89 = {gMainzidev[99:0], 7'h59};
  zdLLziMainzidev8  zdLLziMainzidev8R89 (gzdLLziMainzidev8R89[106:7], gzdLLziMainzidev8R89[6:0], callResR289);
  assign gzdLLziMainzidev8R90 = {gMainzidev[99:0], 7'h5a};
  zdLLziMainzidev8  zdLLziMainzidev8R90 (gzdLLziMainzidev8R90[106:7], gzdLLziMainzidev8R90[6:0], callResR290);
  assign gzdLLziMainzidev8R91 = {gMainzidev[99:0], 7'h5b};
  zdLLziMainzidev8  zdLLziMainzidev8R91 (gzdLLziMainzidev8R91[106:7], gzdLLziMainzidev8R91[6:0], callResR291);
  assign gzdLLziMainzidev8R92 = {gMainzidev[99:0], 7'h5c};
  zdLLziMainzidev8  zdLLziMainzidev8R92 (gzdLLziMainzidev8R92[106:7], gzdLLziMainzidev8R92[6:0], callResR292);
  assign gzdLLziMainzidev8R93 = {gMainzidev[99:0], 7'h5d};
  zdLLziMainzidev8  zdLLziMainzidev8R93 (gzdLLziMainzidev8R93[106:7], gzdLLziMainzidev8R93[6:0], callResR293);
  assign gzdLLziMainzidev8R94 = {gMainzidev[99:0], 7'h5e};
  zdLLziMainzidev8  zdLLziMainzidev8R94 (gzdLLziMainzidev8R94[106:7], gzdLLziMainzidev8R94[6:0], callResR294);
  assign gzdLLziMainzidev8R95 = {gMainzidev[99:0], 7'h5f};
  zdLLziMainzidev8  zdLLziMainzidev8R95 (gzdLLziMainzidev8R95[106:7], gzdLLziMainzidev8R95[6:0], callResR295);
  assign gzdLLziMainzidev8R96 = {gMainzidev[99:0], 7'h60};
  zdLLziMainzidev8  zdLLziMainzidev8R96 (gzdLLziMainzidev8R96[106:7], gzdLLziMainzidev8R96[6:0], callResR296);
  assign gzdLLziMainzidev8R97 = {gMainzidev[99:0], 7'h61};
  zdLLziMainzidev8  zdLLziMainzidev8R97 (gzdLLziMainzidev8R97[106:7], gzdLLziMainzidev8R97[6:0], callResR297);
  assign gzdLLziMainzidev8R98 = {gMainzidev[99:0], 7'h62};
  zdLLziMainzidev8  zdLLziMainzidev8R98 (gzdLLziMainzidev8R98[106:7], gzdLLziMainzidev8R98[6:0], callResR298);
  assign gzdLLziMainzidev8R99 = {gMainzidev[99:0], 7'h63};
  zdLLziMainzidev8  zdLLziMainzidev8R99 (gzdLLziMainzidev8R99[106:7], gzdLLziMainzidev8R99[6:0], callResR299);
  assign gzdLLziMainzidev11 = {gMainzidev[99:0], 7'h00};
  zdLLziMainzidev11  zdLLziMainzidev11 (gzdLLziMainzidev11[106:7], gzdLLziMainzidev11[6:0], callResR300);
  assign gzdLLziMainzidev11R1 = {gMainzidev[99:0], 7'h01};
  zdLLziMainzidev11  zdLLziMainzidev11R1 (gzdLLziMainzidev11R1[106:7], gzdLLziMainzidev11R1[6:0], callResR301);
  assign gzdLLziMainzidev11R2 = {gMainzidev[99:0], 7'h02};
  zdLLziMainzidev11  zdLLziMainzidev11R2 (gzdLLziMainzidev11R2[106:7], gzdLLziMainzidev11R2[6:0], callResR302);
  assign gzdLLziMainzidev11R3 = {gMainzidev[99:0], 7'h03};
  zdLLziMainzidev11  zdLLziMainzidev11R3 (gzdLLziMainzidev11R3[106:7], gzdLLziMainzidev11R3[6:0], callResR303);
  assign gzdLLziMainzidev11R4 = {gMainzidev[99:0], 7'h04};
  zdLLziMainzidev11  zdLLziMainzidev11R4 (gzdLLziMainzidev11R4[106:7], gzdLLziMainzidev11R4[6:0], callResR304);
  assign gzdLLziMainzidev11R5 = {gMainzidev[99:0], 7'h05};
  zdLLziMainzidev11  zdLLziMainzidev11R5 (gzdLLziMainzidev11R5[106:7], gzdLLziMainzidev11R5[6:0], callResR305);
  assign gzdLLziMainzidev11R6 = {gMainzidev[99:0], 7'h06};
  zdLLziMainzidev11  zdLLziMainzidev11R6 (gzdLLziMainzidev11R6[106:7], gzdLLziMainzidev11R6[6:0], callResR306);
  assign gzdLLziMainzidev11R7 = {gMainzidev[99:0], 7'h07};
  zdLLziMainzidev11  zdLLziMainzidev11R7 (gzdLLziMainzidev11R7[106:7], gzdLLziMainzidev11R7[6:0], callResR307);
  assign gzdLLziMainzidev11R8 = {gMainzidev[99:0], 7'h08};
  zdLLziMainzidev11  zdLLziMainzidev11R8 (gzdLLziMainzidev11R8[106:7], gzdLLziMainzidev11R8[6:0], callResR308);
  assign gzdLLziMainzidev11R9 = {gMainzidev[99:0], 7'h09};
  zdLLziMainzidev11  zdLLziMainzidev11R9 (gzdLLziMainzidev11R9[106:7], gzdLLziMainzidev11R9[6:0], callResR309);
  assign gzdLLziMainzidev11R10 = {gMainzidev[99:0], 7'h0a};
  zdLLziMainzidev11  zdLLziMainzidev11R10 (gzdLLziMainzidev11R10[106:7], gzdLLziMainzidev11R10[6:0], callResR310);
  assign gzdLLziMainzidev11R11 = {gMainzidev[99:0], 7'h0b};
  zdLLziMainzidev11  zdLLziMainzidev11R11 (gzdLLziMainzidev11R11[106:7], gzdLLziMainzidev11R11[6:0], callResR311);
  assign gzdLLziMainzidev11R12 = {gMainzidev[99:0], 7'h0c};
  zdLLziMainzidev11  zdLLziMainzidev11R12 (gzdLLziMainzidev11R12[106:7], gzdLLziMainzidev11R12[6:0], callResR312);
  assign gzdLLziMainzidev11R13 = {gMainzidev[99:0], 7'h0d};
  zdLLziMainzidev11  zdLLziMainzidev11R13 (gzdLLziMainzidev11R13[106:7], gzdLLziMainzidev11R13[6:0], callResR313);
  assign gzdLLziMainzidev11R14 = {gMainzidev[99:0], 7'h0e};
  zdLLziMainzidev11  zdLLziMainzidev11R14 (gzdLLziMainzidev11R14[106:7], gzdLLziMainzidev11R14[6:0], callResR314);
  assign gzdLLziMainzidev11R15 = {gMainzidev[99:0], 7'h0f};
  zdLLziMainzidev11  zdLLziMainzidev11R15 (gzdLLziMainzidev11R15[106:7], gzdLLziMainzidev11R15[6:0], callResR315);
  assign gzdLLziMainzidev11R16 = {gMainzidev[99:0], 7'h10};
  zdLLziMainzidev11  zdLLziMainzidev11R16 (gzdLLziMainzidev11R16[106:7], gzdLLziMainzidev11R16[6:0], callResR316);
  assign gzdLLziMainzidev11R17 = {gMainzidev[99:0], 7'h11};
  zdLLziMainzidev11  zdLLziMainzidev11R17 (gzdLLziMainzidev11R17[106:7], gzdLLziMainzidev11R17[6:0], callResR317);
  assign gzdLLziMainzidev11R18 = {gMainzidev[99:0], 7'h12};
  zdLLziMainzidev11  zdLLziMainzidev11R18 (gzdLLziMainzidev11R18[106:7], gzdLLziMainzidev11R18[6:0], callResR318);
  assign gzdLLziMainzidev11R19 = {gMainzidev[99:0], 7'h13};
  zdLLziMainzidev11  zdLLziMainzidev11R19 (gzdLLziMainzidev11R19[106:7], gzdLLziMainzidev11R19[6:0], callResR319);
  assign gzdLLziMainzidev11R20 = {gMainzidev[99:0], 7'h14};
  zdLLziMainzidev11  zdLLziMainzidev11R20 (gzdLLziMainzidev11R20[106:7], gzdLLziMainzidev11R20[6:0], callResR320);
  assign gzdLLziMainzidev11R21 = {gMainzidev[99:0], 7'h15};
  zdLLziMainzidev11  zdLLziMainzidev11R21 (gzdLLziMainzidev11R21[106:7], gzdLLziMainzidev11R21[6:0], callResR321);
  assign gzdLLziMainzidev11R22 = {gMainzidev[99:0], 7'h16};
  zdLLziMainzidev11  zdLLziMainzidev11R22 (gzdLLziMainzidev11R22[106:7], gzdLLziMainzidev11R22[6:0], callResR322);
  assign gzdLLziMainzidev11R23 = {gMainzidev[99:0], 7'h17};
  zdLLziMainzidev11  zdLLziMainzidev11R23 (gzdLLziMainzidev11R23[106:7], gzdLLziMainzidev11R23[6:0], callResR323);
  assign gzdLLziMainzidev11R24 = {gMainzidev[99:0], 7'h18};
  zdLLziMainzidev11  zdLLziMainzidev11R24 (gzdLLziMainzidev11R24[106:7], gzdLLziMainzidev11R24[6:0], callResR324);
  assign gzdLLziMainzidev11R25 = {gMainzidev[99:0], 7'h19};
  zdLLziMainzidev11  zdLLziMainzidev11R25 (gzdLLziMainzidev11R25[106:7], gzdLLziMainzidev11R25[6:0], callResR325);
  assign gzdLLziMainzidev11R26 = {gMainzidev[99:0], 7'h1a};
  zdLLziMainzidev11  zdLLziMainzidev11R26 (gzdLLziMainzidev11R26[106:7], gzdLLziMainzidev11R26[6:0], callResR326);
  assign gzdLLziMainzidev11R27 = {gMainzidev[99:0], 7'h1b};
  zdLLziMainzidev11  zdLLziMainzidev11R27 (gzdLLziMainzidev11R27[106:7], gzdLLziMainzidev11R27[6:0], callResR327);
  assign gzdLLziMainzidev11R28 = {gMainzidev[99:0], 7'h1c};
  zdLLziMainzidev11  zdLLziMainzidev11R28 (gzdLLziMainzidev11R28[106:7], gzdLLziMainzidev11R28[6:0], callResR328);
  assign gzdLLziMainzidev11R29 = {gMainzidev[99:0], 7'h1d};
  zdLLziMainzidev11  zdLLziMainzidev11R29 (gzdLLziMainzidev11R29[106:7], gzdLLziMainzidev11R29[6:0], callResR329);
  assign gzdLLziMainzidev11R30 = {gMainzidev[99:0], 7'h1e};
  zdLLziMainzidev11  zdLLziMainzidev11R30 (gzdLLziMainzidev11R30[106:7], gzdLLziMainzidev11R30[6:0], callResR330);
  assign gzdLLziMainzidev11R31 = {gMainzidev[99:0], 7'h1f};
  zdLLziMainzidev11  zdLLziMainzidev11R31 (gzdLLziMainzidev11R31[106:7], gzdLLziMainzidev11R31[6:0], callResR331);
  assign gzdLLziMainzidev11R32 = {gMainzidev[99:0], 7'h20};
  zdLLziMainzidev11  zdLLziMainzidev11R32 (gzdLLziMainzidev11R32[106:7], gzdLLziMainzidev11R32[6:0], callResR332);
  assign gzdLLziMainzidev11R33 = {gMainzidev[99:0], 7'h21};
  zdLLziMainzidev11  zdLLziMainzidev11R33 (gzdLLziMainzidev11R33[106:7], gzdLLziMainzidev11R33[6:0], callResR333);
  assign gzdLLziMainzidev11R34 = {gMainzidev[99:0], 7'h22};
  zdLLziMainzidev11  zdLLziMainzidev11R34 (gzdLLziMainzidev11R34[106:7], gzdLLziMainzidev11R34[6:0], callResR334);
  assign gzdLLziMainzidev11R35 = {gMainzidev[99:0], 7'h23};
  zdLLziMainzidev11  zdLLziMainzidev11R35 (gzdLLziMainzidev11R35[106:7], gzdLLziMainzidev11R35[6:0], callResR335);
  assign gzdLLziMainzidev11R36 = {gMainzidev[99:0], 7'h24};
  zdLLziMainzidev11  zdLLziMainzidev11R36 (gzdLLziMainzidev11R36[106:7], gzdLLziMainzidev11R36[6:0], callResR336);
  assign gzdLLziMainzidev11R37 = {gMainzidev[99:0], 7'h25};
  zdLLziMainzidev11  zdLLziMainzidev11R37 (gzdLLziMainzidev11R37[106:7], gzdLLziMainzidev11R37[6:0], callResR337);
  assign gzdLLziMainzidev11R38 = {gMainzidev[99:0], 7'h26};
  zdLLziMainzidev11  zdLLziMainzidev11R38 (gzdLLziMainzidev11R38[106:7], gzdLLziMainzidev11R38[6:0], callResR338);
  assign gzdLLziMainzidev11R39 = {gMainzidev[99:0], 7'h27};
  zdLLziMainzidev11  zdLLziMainzidev11R39 (gzdLLziMainzidev11R39[106:7], gzdLLziMainzidev11R39[6:0], callResR339);
  assign gzdLLziMainzidev11R40 = {gMainzidev[99:0], 7'h28};
  zdLLziMainzidev11  zdLLziMainzidev11R40 (gzdLLziMainzidev11R40[106:7], gzdLLziMainzidev11R40[6:0], callResR340);
  assign gzdLLziMainzidev11R41 = {gMainzidev[99:0], 7'h29};
  zdLLziMainzidev11  zdLLziMainzidev11R41 (gzdLLziMainzidev11R41[106:7], gzdLLziMainzidev11R41[6:0], callResR341);
  assign gzdLLziMainzidev11R42 = {gMainzidev[99:0], 7'h2a};
  zdLLziMainzidev11  zdLLziMainzidev11R42 (gzdLLziMainzidev11R42[106:7], gzdLLziMainzidev11R42[6:0], callResR342);
  assign gzdLLziMainzidev11R43 = {gMainzidev[99:0], 7'h2b};
  zdLLziMainzidev11  zdLLziMainzidev11R43 (gzdLLziMainzidev11R43[106:7], gzdLLziMainzidev11R43[6:0], callResR343);
  assign gzdLLziMainzidev11R44 = {gMainzidev[99:0], 7'h2c};
  zdLLziMainzidev11  zdLLziMainzidev11R44 (gzdLLziMainzidev11R44[106:7], gzdLLziMainzidev11R44[6:0], callResR344);
  assign gzdLLziMainzidev11R45 = {gMainzidev[99:0], 7'h2d};
  zdLLziMainzidev11  zdLLziMainzidev11R45 (gzdLLziMainzidev11R45[106:7], gzdLLziMainzidev11R45[6:0], callResR345);
  assign gzdLLziMainzidev11R46 = {gMainzidev[99:0], 7'h2e};
  zdLLziMainzidev11  zdLLziMainzidev11R46 (gzdLLziMainzidev11R46[106:7], gzdLLziMainzidev11R46[6:0], callResR346);
  assign gzdLLziMainzidev11R47 = {gMainzidev[99:0], 7'h2f};
  zdLLziMainzidev11  zdLLziMainzidev11R47 (gzdLLziMainzidev11R47[106:7], gzdLLziMainzidev11R47[6:0], callResR347);
  assign gzdLLziMainzidev11R48 = {gMainzidev[99:0], 7'h30};
  zdLLziMainzidev11  zdLLziMainzidev11R48 (gzdLLziMainzidev11R48[106:7], gzdLLziMainzidev11R48[6:0], callResR348);
  assign gzdLLziMainzidev11R49 = {gMainzidev[99:0], 7'h31};
  zdLLziMainzidev11  zdLLziMainzidev11R49 (gzdLLziMainzidev11R49[106:7], gzdLLziMainzidev11R49[6:0], callResR349);
  assign gzdLLziMainzidev11R50 = {gMainzidev[99:0], 7'h32};
  zdLLziMainzidev11  zdLLziMainzidev11R50 (gzdLLziMainzidev11R50[106:7], gzdLLziMainzidev11R50[6:0], callResR350);
  assign gzdLLziMainzidev11R51 = {gMainzidev[99:0], 7'h33};
  zdLLziMainzidev11  zdLLziMainzidev11R51 (gzdLLziMainzidev11R51[106:7], gzdLLziMainzidev11R51[6:0], callResR351);
  assign gzdLLziMainzidev11R52 = {gMainzidev[99:0], 7'h34};
  zdLLziMainzidev11  zdLLziMainzidev11R52 (gzdLLziMainzidev11R52[106:7], gzdLLziMainzidev11R52[6:0], callResR352);
  assign gzdLLziMainzidev11R53 = {gMainzidev[99:0], 7'h35};
  zdLLziMainzidev11  zdLLziMainzidev11R53 (gzdLLziMainzidev11R53[106:7], gzdLLziMainzidev11R53[6:0], callResR353);
  assign gzdLLziMainzidev11R54 = {gMainzidev[99:0], 7'h36};
  zdLLziMainzidev11  zdLLziMainzidev11R54 (gzdLLziMainzidev11R54[106:7], gzdLLziMainzidev11R54[6:0], callResR354);
  assign gzdLLziMainzidev11R55 = {gMainzidev[99:0], 7'h37};
  zdLLziMainzidev11  zdLLziMainzidev11R55 (gzdLLziMainzidev11R55[106:7], gzdLLziMainzidev11R55[6:0], callResR355);
  assign gzdLLziMainzidev11R56 = {gMainzidev[99:0], 7'h38};
  zdLLziMainzidev11  zdLLziMainzidev11R56 (gzdLLziMainzidev11R56[106:7], gzdLLziMainzidev11R56[6:0], callResR356);
  assign gzdLLziMainzidev11R57 = {gMainzidev[99:0], 7'h39};
  zdLLziMainzidev11  zdLLziMainzidev11R57 (gzdLLziMainzidev11R57[106:7], gzdLLziMainzidev11R57[6:0], callResR357);
  assign gzdLLziMainzidev11R58 = {gMainzidev[99:0], 7'h3a};
  zdLLziMainzidev11  zdLLziMainzidev11R58 (gzdLLziMainzidev11R58[106:7], gzdLLziMainzidev11R58[6:0], callResR358);
  assign gzdLLziMainzidev11R59 = {gMainzidev[99:0], 7'h3b};
  zdLLziMainzidev11  zdLLziMainzidev11R59 (gzdLLziMainzidev11R59[106:7], gzdLLziMainzidev11R59[6:0], callResR359);
  assign gzdLLziMainzidev11R60 = {gMainzidev[99:0], 7'h3c};
  zdLLziMainzidev11  zdLLziMainzidev11R60 (gzdLLziMainzidev11R60[106:7], gzdLLziMainzidev11R60[6:0], callResR360);
  assign gzdLLziMainzidev11R61 = {gMainzidev[99:0], 7'h3d};
  zdLLziMainzidev11  zdLLziMainzidev11R61 (gzdLLziMainzidev11R61[106:7], gzdLLziMainzidev11R61[6:0], callResR361);
  assign gzdLLziMainzidev11R62 = {gMainzidev[99:0], 7'h3e};
  zdLLziMainzidev11  zdLLziMainzidev11R62 (gzdLLziMainzidev11R62[106:7], gzdLLziMainzidev11R62[6:0], callResR362);
  assign gzdLLziMainzidev11R63 = {gMainzidev[99:0], 7'h3f};
  zdLLziMainzidev11  zdLLziMainzidev11R63 (gzdLLziMainzidev11R63[106:7], gzdLLziMainzidev11R63[6:0], callResR363);
  assign gzdLLziMainzidev11R64 = {gMainzidev[99:0], 7'h40};
  zdLLziMainzidev11  zdLLziMainzidev11R64 (gzdLLziMainzidev11R64[106:7], gzdLLziMainzidev11R64[6:0], callResR364);
  assign gzdLLziMainzidev11R65 = {gMainzidev[99:0], 7'h41};
  zdLLziMainzidev11  zdLLziMainzidev11R65 (gzdLLziMainzidev11R65[106:7], gzdLLziMainzidev11R65[6:0], callResR365);
  assign gzdLLziMainzidev11R66 = {gMainzidev[99:0], 7'h42};
  zdLLziMainzidev11  zdLLziMainzidev11R66 (gzdLLziMainzidev11R66[106:7], gzdLLziMainzidev11R66[6:0], callResR366);
  assign gzdLLziMainzidev11R67 = {gMainzidev[99:0], 7'h43};
  zdLLziMainzidev11  zdLLziMainzidev11R67 (gzdLLziMainzidev11R67[106:7], gzdLLziMainzidev11R67[6:0], callResR367);
  assign gzdLLziMainzidev11R68 = {gMainzidev[99:0], 7'h44};
  zdLLziMainzidev11  zdLLziMainzidev11R68 (gzdLLziMainzidev11R68[106:7], gzdLLziMainzidev11R68[6:0], callResR368);
  assign gzdLLziMainzidev11R69 = {gMainzidev[99:0], 7'h45};
  zdLLziMainzidev11  zdLLziMainzidev11R69 (gzdLLziMainzidev11R69[106:7], gzdLLziMainzidev11R69[6:0], callResR369);
  assign gzdLLziMainzidev11R70 = {gMainzidev[99:0], 7'h46};
  zdLLziMainzidev11  zdLLziMainzidev11R70 (gzdLLziMainzidev11R70[106:7], gzdLLziMainzidev11R70[6:0], callResR370);
  assign gzdLLziMainzidev11R71 = {gMainzidev[99:0], 7'h47};
  zdLLziMainzidev11  zdLLziMainzidev11R71 (gzdLLziMainzidev11R71[106:7], gzdLLziMainzidev11R71[6:0], callResR371);
  assign gzdLLziMainzidev11R72 = {gMainzidev[99:0], 7'h48};
  zdLLziMainzidev11  zdLLziMainzidev11R72 (gzdLLziMainzidev11R72[106:7], gzdLLziMainzidev11R72[6:0], callResR372);
  assign gzdLLziMainzidev11R73 = {gMainzidev[99:0], 7'h49};
  zdLLziMainzidev11  zdLLziMainzidev11R73 (gzdLLziMainzidev11R73[106:7], gzdLLziMainzidev11R73[6:0], callResR373);
  assign gzdLLziMainzidev11R74 = {gMainzidev[99:0], 7'h4a};
  zdLLziMainzidev11  zdLLziMainzidev11R74 (gzdLLziMainzidev11R74[106:7], gzdLLziMainzidev11R74[6:0], callResR374);
  assign gzdLLziMainzidev11R75 = {gMainzidev[99:0], 7'h4b};
  zdLLziMainzidev11  zdLLziMainzidev11R75 (gzdLLziMainzidev11R75[106:7], gzdLLziMainzidev11R75[6:0], callResR375);
  assign gzdLLziMainzidev11R76 = {gMainzidev[99:0], 7'h4c};
  zdLLziMainzidev11  zdLLziMainzidev11R76 (gzdLLziMainzidev11R76[106:7], gzdLLziMainzidev11R76[6:0], callResR376);
  assign gzdLLziMainzidev11R77 = {gMainzidev[99:0], 7'h4d};
  zdLLziMainzidev11  zdLLziMainzidev11R77 (gzdLLziMainzidev11R77[106:7], gzdLLziMainzidev11R77[6:0], callResR377);
  assign gzdLLziMainzidev11R78 = {gMainzidev[99:0], 7'h4e};
  zdLLziMainzidev11  zdLLziMainzidev11R78 (gzdLLziMainzidev11R78[106:7], gzdLLziMainzidev11R78[6:0], callResR378);
  assign gzdLLziMainzidev11R79 = {gMainzidev[99:0], 7'h4f};
  zdLLziMainzidev11  zdLLziMainzidev11R79 (gzdLLziMainzidev11R79[106:7], gzdLLziMainzidev11R79[6:0], callResR379);
  assign gzdLLziMainzidev11R80 = {gMainzidev[99:0], 7'h50};
  zdLLziMainzidev11  zdLLziMainzidev11R80 (gzdLLziMainzidev11R80[106:7], gzdLLziMainzidev11R80[6:0], callResR380);
  assign gzdLLziMainzidev11R81 = {gMainzidev[99:0], 7'h51};
  zdLLziMainzidev11  zdLLziMainzidev11R81 (gzdLLziMainzidev11R81[106:7], gzdLLziMainzidev11R81[6:0], callResR381);
  assign gzdLLziMainzidev11R82 = {gMainzidev[99:0], 7'h52};
  zdLLziMainzidev11  zdLLziMainzidev11R82 (gzdLLziMainzidev11R82[106:7], gzdLLziMainzidev11R82[6:0], callResR382);
  assign gzdLLziMainzidev11R83 = {gMainzidev[99:0], 7'h53};
  zdLLziMainzidev11  zdLLziMainzidev11R83 (gzdLLziMainzidev11R83[106:7], gzdLLziMainzidev11R83[6:0], callResR383);
  assign gzdLLziMainzidev11R84 = {gMainzidev[99:0], 7'h54};
  zdLLziMainzidev11  zdLLziMainzidev11R84 (gzdLLziMainzidev11R84[106:7], gzdLLziMainzidev11R84[6:0], callResR384);
  assign gzdLLziMainzidev11R85 = {gMainzidev[99:0], 7'h55};
  zdLLziMainzidev11  zdLLziMainzidev11R85 (gzdLLziMainzidev11R85[106:7], gzdLLziMainzidev11R85[6:0], callResR385);
  assign gzdLLziMainzidev11R86 = {gMainzidev[99:0], 7'h56};
  zdLLziMainzidev11  zdLLziMainzidev11R86 (gzdLLziMainzidev11R86[106:7], gzdLLziMainzidev11R86[6:0], callResR386);
  assign gzdLLziMainzidev11R87 = {gMainzidev[99:0], 7'h57};
  zdLLziMainzidev11  zdLLziMainzidev11R87 (gzdLLziMainzidev11R87[106:7], gzdLLziMainzidev11R87[6:0], callResR387);
  assign gzdLLziMainzidev11R88 = {gMainzidev[99:0], 7'h58};
  zdLLziMainzidev11  zdLLziMainzidev11R88 (gzdLLziMainzidev11R88[106:7], gzdLLziMainzidev11R88[6:0], callResR388);
  assign gzdLLziMainzidev11R89 = {gMainzidev[99:0], 7'h59};
  zdLLziMainzidev11  zdLLziMainzidev11R89 (gzdLLziMainzidev11R89[106:7], gzdLLziMainzidev11R89[6:0], callResR389);
  assign gzdLLziMainzidev11R90 = {gMainzidev[99:0], 7'h5a};
  zdLLziMainzidev11  zdLLziMainzidev11R90 (gzdLLziMainzidev11R90[106:7], gzdLLziMainzidev11R90[6:0], callResR390);
  assign gzdLLziMainzidev11R91 = {gMainzidev[99:0], 7'h5b};
  zdLLziMainzidev11  zdLLziMainzidev11R91 (gzdLLziMainzidev11R91[106:7], gzdLLziMainzidev11R91[6:0], callResR391);
  assign gzdLLziMainzidev11R92 = {gMainzidev[99:0], 7'h5c};
  zdLLziMainzidev11  zdLLziMainzidev11R92 (gzdLLziMainzidev11R92[106:7], gzdLLziMainzidev11R92[6:0], callResR392);
  assign gzdLLziMainzidev11R93 = {gMainzidev[99:0], 7'h5d};
  zdLLziMainzidev11  zdLLziMainzidev11R93 (gzdLLziMainzidev11R93[106:7], gzdLLziMainzidev11R93[6:0], callResR393);
  assign gzdLLziMainzidev11R94 = {gMainzidev[99:0], 7'h5e};
  zdLLziMainzidev11  zdLLziMainzidev11R94 (gzdLLziMainzidev11R94[106:7], gzdLLziMainzidev11R94[6:0], callResR394);
  assign gzdLLziMainzidev11R95 = {gMainzidev[99:0], 7'h5f};
  zdLLziMainzidev11  zdLLziMainzidev11R95 (gzdLLziMainzidev11R95[106:7], gzdLLziMainzidev11R95[6:0], callResR395);
  assign gzdLLziMainzidev11R96 = {gMainzidev[99:0], 7'h60};
  zdLLziMainzidev11  zdLLziMainzidev11R96 (gzdLLziMainzidev11R96[106:7], gzdLLziMainzidev11R96[6:0], callResR396);
  assign gzdLLziMainzidev11R97 = {gMainzidev[99:0], 7'h61};
  zdLLziMainzidev11  zdLLziMainzidev11R97 (gzdLLziMainzidev11R97[106:7], gzdLLziMainzidev11R97[6:0], callResR397);
  assign gzdLLziMainzidev11R98 = {gMainzidev[99:0], 7'h62};
  zdLLziMainzidev11  zdLLziMainzidev11R98 (gzdLLziMainzidev11R98[106:7], gzdLLziMainzidev11R98[6:0], callResR398);
  assign gzdLLziMainzidev11R99 = {gMainzidev[99:0], 7'h63};
  zdLLziMainzidev11  zdLLziMainzidev11R99 (gzdLLziMainzidev11R99[106:7], gzdLLziMainzidev11R99[6:0], callResR399);
  assign {__continue, __out0, __out1, __out2, __out3, __resumption_tag_next} = {1'h1, callRes, callResR1, callResR2, callResR3, callResR4, callResR5, callResR6, callResR7, callResR8, callResR9, callResR10, callResR11, callResR12, callResR13, callResR14, callResR15, callResR16, callResR17, callResR18, callResR19, callResR20, callResR21, callResR22, callResR23, callResR24, callResR25, callResR26, callResR27, callResR28, callResR29, callResR30, callResR31, callResR32, callResR33, callResR34, callResR35, callResR36, callResR37, callResR38, callResR39, callResR40, callResR41, callResR42, callResR43, callResR44, callResR45, callResR46, callResR47, callResR48, callResR49, callResR50, callResR51, callResR52, callResR53, callResR54, callResR55, callResR56, callResR57, callResR58, callResR59, callResR60, callResR61, callResR62, callResR63, callResR64, callResR65, callResR66, callResR67, callResR68, callResR69, callResR70, callResR71, callResR72, callResR73, callResR74, callResR75, callResR76, callResR77, callResR78, callResR79, callResR80, callResR81, callResR82, callResR83, callResR84, callResR85, callResR86, callResR87, callResR88, callResR89, callResR90, callResR91, callResR92, callResR93, callResR94, callResR95, callResR96, callResR97, callResR98, callResR99, callResR100, callResR101, callResR102, callResR103, callResR104, callResR105, callResR106, callResR107, callResR108, callResR109, callResR110, callResR111, callResR112, callResR113, callResR114, callResR115, callResR116, callResR117, callResR118, callResR119, callResR120, callResR121, callResR122, callResR123, callResR124, callResR125, callResR126, callResR127, callResR128, callResR129, callResR130, callResR131, callResR132, callResR133, callResR134, callResR135, callResR136, callResR137, callResR138, callResR139, callResR140, callResR141, callResR142, callResR143, callResR144, callResR145, callResR146, callResR147, callResR148, callResR149, callResR150, callResR151, callResR152, callResR153, callResR154, callResR155, callResR156, callResR157, callResR158, callResR159, callResR160, callResR161, callResR162, callResR163, callResR164, callResR165, callResR166, callResR167, callResR168, callResR169, callResR170, callResR171, callResR172, callResR173, callResR174, callResR175, callResR176, callResR177, callResR178, callResR179, callResR180, callResR181, callResR182, callResR183, callResR184, callResR185, callResR186, callResR187, callResR188, callResR189, callResR190, callResR191, callResR192, callResR193, callResR194, callResR195, callResR196, callResR197, callResR198, callResR199, callResR200, callResR201, callResR202, callResR203, callResR204, callResR205, callResR206, callResR207, callResR208, callResR209, callResR210, callResR211, callResR212, callResR213, callResR214, callResR215, callResR216, callResR217, callResR218, callResR219, callResR220, callResR221, callResR222, callResR223, callResR224, callResR225, callResR226, callResR227, callResR228, callResR229, callResR230, callResR231, callResR232, callResR233, callResR234, callResR235, callResR236, callResR237, callResR238, callResR239, callResR240, callResR241, callResR242, callResR243, callResR244, callResR245, callResR246, callResR247, callResR248, callResR249, callResR250, callResR251, callResR252, callResR253, callResR254, callResR255, callResR256, callResR257, callResR258, callResR259, callResR260, callResR261, callResR262, callResR263, callResR264, callResR265, callResR266, callResR267, callResR268, callResR269, callResR270, callResR271, callResR272, callResR273, callResR274, callResR275, callResR276, callResR277, callResR278, callResR279, callResR280, callResR281, callResR282, callResR283, callResR284, callResR285, callResR286, callResR287, callResR288, callResR289, callResR290, callResR291, callResR292, callResR293, callResR294, callResR295, callResR296, callResR297, callResR298, callResR299, callResR300, callResR301, callResR302, callResR303, callResR304, callResR305, callResR306, callResR307, callResR308, callResR309, callResR310, callResR311, callResR312, callResR313, callResR314, callResR315, callResR316, callResR317, callResR318, callResR319, callResR320, callResR321, callResR322, callResR323, callResR324, callResR325, callResR326, callResR327, callResR328, callResR329, callResR330, callResR331, callResR332, callResR333, callResR334, callResR335, callResR336, callResR337, callResR338, callResR339, callResR340, callResR341, callResR342, callResR343, callResR344, callResR345, callResR346, callResR347, callResR348, callResR349, callResR350, callResR351, callResR352, callResR353, callResR354, callResR355, callResR356, callResR357, callResR358, callResR359, callResR360, callResR361, callResR362, callResR363, callResR364, callResR365, callResR366, callResR367, callResR368, callResR369, callResR370, callResR371, callResR372, callResR373, callResR374, callResR375, callResR376, callResR377, callResR378, callResR379, callResR380, callResR381, callResR382, callResR383, callResR384, callResR385, callResR386, callResR387, callResR388, callResR389, callResR390, callResR391, callResR392, callResR393, callResR394, callResR395, callResR396, callResR397, callResR398, callResR399};
  initial __resumption_tag <= {7'h64{1'h0}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      __resumption_tag <= {7'h64{1'h0}};
    end else begin
      __resumption_tag <= __resumption_tag_next;
    end
  end
endmodule

module zdLLziMainzidev2 (input logic [99:0] arg0,
  input logic [6:0] arg1,
  output logic [0:0] res);
  logic [6:0] resizze;
  logic [127:0] resizzeR1;
  logic [0:0] msbit;
  logic [0:0] gReWireziPreludezinot;
  logic [0:0] callRes;
  logic [6:0] resizzeR2;
  logic [127:0] resizzeR3;
  logic [0:0] msbitR1;
  logic [0:0] gReWireziPreludezinotR1;
  logic [0:0] callResR1;
  logic [107:0] gzdLLziMainzidev1;
  logic [99:0] gMainzix2;
  logic [99:0] callResR2;
  logic [99:0] resizzeR4;
  logic [6:0] resizzeR5;
  logic [255:0] binOp;
  logic [255:0] binOpR1;
  logic [127:0] resizzeR6;
  logic [6:0] resizzeR7;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR8;
  logic [6:0] resizzeR9;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [127:0] resizzeR10;
  logic [107:0] gzdLLziMainzidev;
  logic [99:0] resizzeR11;
  logic [6:0] resizzeR12;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [127:0] resizzeR13;
  logic [6:0] resizzeR14;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [127:0] resizzeR15;
  assign resizze = arg1;
  assign resizzeR1 = 128'(resizze[6:0]);
  assign msbit = resizzeR1[0];
  assign gReWireziPreludezinot = msbit[0];
  ReWireziPreludezinot  ReWireziPreludezinot (gReWireziPreludezinot[0], callRes);
  assign resizzeR2 = arg1;
  assign resizzeR3 = 128'(resizzeR2[6:0]);
  assign msbitR1 = resizzeR3[0];
  assign gReWireziPreludezinotR1 = msbitR1[0];
  ReWireziPreludezinot  ReWireziPreludezinotR1 (gReWireziPreludezinotR1[0], callResR1);
  assign gzdLLziMainzidev1 = {arg0, arg1, callResR1};
  assign gMainzix2 = gzdLLziMainzidev1[107:8];
  Mainzix2  Mainzix2 (gMainzix2[99:0], callResR2);
  assign resizzeR4 = callResR2;
  assign resizzeR5 = gzdLLziMainzidev1[7:1];
  assign binOp = {128'(resizzeR5[6:0]), 128'h00000000000000000000000000000001};
  assign binOpR1 = {binOp[255:128] - binOp[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR6 = binOpR1[255:128] % binOpR1[127:0];
  assign resizzeR7 = resizzeR6[6:0];
  assign binOpR2 = {128'(resizzeR7[6:0]), 128'h00000000000000000000000000000002};
  assign binOpR3 = {binOpR2[255:128] / binOpR2[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR8 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR9 = resizzeR8[6:0];
  assign binOpR4 = {128'h00000000000000000000000000000064, 128'(resizzeR9[6:0])};
  assign binOpR5 = {binOpR4[255:128] - binOpR4[127:0], 128'h00000000000000000000000000000001};
  assign binOpR6 = {binOpR5[255:128] - binOpR5[127:0], 128'h00000000000000000000000000000001};
  assign binOpR7 = {128'(resizzeR4[99:0]), binOpR6[255:128] * binOpR6[127:0]};
  assign resizzeR10 = binOpR7[255:128] >> binOpR7[127:0];
  assign gzdLLziMainzidev = {arg0, arg1, callRes};
  assign resizzeR11 = gzdLLziMainzidev[107:8];
  assign resizzeR12 = gzdLLziMainzidev[7:1];
  assign binOpR8 = {128'(resizzeR12[6:0]), 128'h00000000000000000000000000000002};
  assign binOpR9 = {binOpR8[255:128] / binOpR8[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR13 = binOpR9[255:128] % binOpR9[127:0];
  assign resizzeR14 = resizzeR13[6:0];
  assign binOpR10 = {128'h00000000000000000000000000000064, 128'(resizzeR14[6:0])};
  assign binOpR11 = {binOpR10[255:128] - binOpR10[127:0], 128'h00000000000000000000000000000001};
  assign binOpR12 = {binOpR11[255:128] - binOpR11[127:0], 128'h00000000000000000000000000000001};
  assign binOpR13 = {128'(resizzeR11[99:0]), binOpR12[255:128] * binOpR12[127:0]};
  assign resizzeR15 = binOpR13[255:128] >> binOpR13[127:0];
  assign res = (gzdLLziMainzidev[0] == 1'h1) ? resizzeR15[0] : resizzeR10[0];
endmodule

module zdLLziMainzidev5 (input logic [99:0] arg0,
  input logic [6:0] arg1,
  output logic [0:0] res);
  logic [6:0] resizze;
  logic [127:0] resizzeR1;
  logic [0:0] msbit;
  logic [0:0] gReWireziPreludezinot;
  logic [0:0] callRes;
  logic [6:0] resizzeR2;
  logic [127:0] resizzeR3;
  logic [0:0] msbitR1;
  logic [0:0] gReWireziPreludezinotR1;
  logic [0:0] callResR1;
  logic [107:0] gzdLLziMainzidev4;
  logic [99:0] gMainzix2;
  logic [99:0] callResR2;
  logic [99:0] resizzeR4;
  logic [6:0] resizzeR5;
  logic [255:0] binOp;
  logic [255:0] binOpR1;
  logic [127:0] resizzeR6;
  logic [6:0] resizzeR7;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR8;
  logic [6:0] resizzeR9;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR10;
  logic [6:0] resizzeR11;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [127:0] resizzeR12;
  logic [107:0] gzdLLziMainzidev3;
  logic [99:0] resizzeR13;
  logic [6:0] resizzeR14;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [127:0] resizzeR15;
  logic [6:0] resizzeR16;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [127:0] resizzeR17;
  logic [6:0] resizzeR18;
  logic [255:0] binOpR14;
  logic [255:0] binOpR15;
  logic [255:0] binOpR16;
  logic [255:0] binOpR17;
  logic [127:0] resizzeR19;
  assign resizze = arg1;
  assign resizzeR1 = 128'(resizze[6:0]);
  assign msbit = resizzeR1[0];
  assign gReWireziPreludezinot = msbit[0];
  ReWireziPreludezinot  ReWireziPreludezinot (gReWireziPreludezinot[0], callRes);
  assign resizzeR2 = arg1;
  assign resizzeR3 = 128'(resizzeR2[6:0]);
  assign msbitR1 = resizzeR3[0];
  assign gReWireziPreludezinotR1 = msbitR1[0];
  ReWireziPreludezinot  ReWireziPreludezinotR1 (gReWireziPreludezinotR1[0], callResR1);
  assign gzdLLziMainzidev4 = {arg0, arg1, callResR1};
  assign gMainzix2 = gzdLLziMainzidev4[107:8];
  Mainzix2  Mainzix2 (gMainzix2[99:0], callResR2);
  assign resizzeR4 = callResR2;
  assign resizzeR5 = gzdLLziMainzidev4[7:1];
  assign binOp = {128'(resizzeR5[6:0]), 128'h00000000000000000000000000000001};
  assign binOpR1 = {binOp[255:128] - binOp[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR6 = binOpR1[255:128] % binOpR1[127:0];
  assign resizzeR7 = resizzeR6[6:0];
  assign binOpR2 = {128'h00000000000000000000000000000031, 128'(resizzeR7[6:0])};
  assign binOpR3 = {binOpR2[255:128] + binOpR2[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR8 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR9 = resizzeR8[6:0];
  assign binOpR4 = {128'(resizzeR9[6:0]), 128'h00000000000000000000000000000002};
  assign binOpR5 = {binOpR4[255:128] / binOpR4[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR10 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR11 = resizzeR10[6:0];
  assign binOpR6 = {128'h00000000000000000000000000000064, 128'(resizzeR11[6:0])};
  assign binOpR7 = {binOpR6[255:128] - binOpR6[127:0], 128'h00000000000000000000000000000001};
  assign binOpR8 = {binOpR7[255:128] - binOpR7[127:0], 128'h00000000000000000000000000000001};
  assign binOpR9 = {128'(resizzeR4[99:0]), binOpR8[255:128] * binOpR8[127:0]};
  assign resizzeR12 = binOpR9[255:128] >> binOpR9[127:0];
  assign gzdLLziMainzidev3 = {arg0, arg1, callRes};
  assign resizzeR13 = gzdLLziMainzidev3[107:8];
  assign resizzeR14 = gzdLLziMainzidev3[7:1];
  assign binOpR10 = {128'h00000000000000000000000000000031, 128'(resizzeR14[6:0])};
  assign binOpR11 = {binOpR10[255:128] + binOpR10[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR15 = binOpR11[255:128] % binOpR11[127:0];
  assign resizzeR16 = resizzeR15[6:0];
  assign binOpR12 = {128'(resizzeR16[6:0]), 128'h00000000000000000000000000000002};
  assign binOpR13 = {binOpR12[255:128] / binOpR12[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR17 = binOpR13[255:128] % binOpR13[127:0];
  assign resizzeR18 = resizzeR17[6:0];
  assign binOpR14 = {128'h00000000000000000000000000000064, 128'(resizzeR18[6:0])};
  assign binOpR15 = {binOpR14[255:128] - binOpR14[127:0], 128'h00000000000000000000000000000001};
  assign binOpR16 = {binOpR15[255:128] - binOpR15[127:0], 128'h00000000000000000000000000000001};
  assign binOpR17 = {128'(resizzeR13[99:0]), binOpR16[255:128] * binOpR16[127:0]};
  assign resizzeR19 = binOpR17[255:128] >> binOpR17[127:0];
  assign res = (gzdLLziMainzidev3[0] == 1'h1) ? resizzeR19[0] : resizzeR12[0];
endmodule

module zdLLziMainzidev8 (input logic [99:0] arg0,
  input logic [6:0] arg1,
  output logic [0:0] res);
  logic [6:0] resizze;
  logic [255:0] binOp;
  logic [6:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [107:0] gzdLLziMainzidev7;
  logic [99:0] gMainzix2;
  logic [99:0] callRes;
  logic [99:0] resizzeR2;
  logic [6:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [6:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR6;
  logic [6:0] resizzeR7;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [127:0] resizzeR8;
  logic [107:0] gzdLLziMainzidev6;
  logic [99:0] resizzeR9;
  logic [6:0] resizzeR10;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [127:0] resizzeR11;
  logic [6:0] resizzeR12;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [255:0] binOpR14;
  logic [255:0] binOpR15;
  logic [127:0] resizzeR13;
  assign resizze = arg1;
  assign binOp = {128'(resizze[6:0]), 128'h00000000000000000000000000000031};
  assign resizzeR1 = arg1;
  assign binOpR1 = {128'(resizzeR1[6:0]), 128'h00000000000000000000000000000031};
  assign gzdLLziMainzidev7 = {arg0, arg1, binOpR1[255:128] < binOpR1[127:0]};
  assign gMainzix2 = gzdLLziMainzidev7[107:8];
  Mainzix2  Mainzix2 (gMainzix2[99:0], callRes);
  assign resizzeR2 = callRes;
  assign resizzeR3 = gzdLLziMainzidev7[7:1];
  assign binOpR2 = {128'(resizzeR3[6:0]), 128'h00000000000000000000000000000031};
  assign binOpR3 = {binOpR2[255:128] - binOpR2[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[6:0];
  assign binOpR4 = {128'(resizzeR5[6:0]), 128'h00000000000000000000000000000002};
  assign binOpR5 = {binOpR4[255:128] * binOpR4[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR6 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR7 = resizzeR6[6:0];
  assign binOpR6 = {128'h00000000000000000000000000000064, 128'(resizzeR7[6:0])};
  assign binOpR7 = {binOpR6[255:128] - binOpR6[127:0], 128'h00000000000000000000000000000001};
  assign binOpR8 = {binOpR7[255:128] - binOpR7[127:0], 128'h00000000000000000000000000000001};
  assign binOpR9 = {128'(resizzeR2[99:0]), binOpR8[255:128] * binOpR8[127:0]};
  assign resizzeR8 = binOpR9[255:128] >> binOpR9[127:0];
  assign gzdLLziMainzidev6 = {arg0, arg1, binOp[255:128] < binOp[127:0]};
  assign resizzeR9 = gzdLLziMainzidev6[107:8];
  assign resizzeR10 = gzdLLziMainzidev6[7:1];
  assign binOpR10 = {128'(resizzeR10[6:0]), 128'h00000000000000000000000000000002};
  assign binOpR11 = {binOpR10[255:128] * binOpR10[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR11 = binOpR11[255:128] % binOpR11[127:0];
  assign resizzeR12 = resizzeR11[6:0];
  assign binOpR12 = {128'h00000000000000000000000000000064, 128'(resizzeR12[6:0])};
  assign binOpR13 = {binOpR12[255:128] - binOpR12[127:0], 128'h00000000000000000000000000000001};
  assign binOpR14 = {binOpR13[255:128] - binOpR13[127:0], 128'h00000000000000000000000000000001};
  assign binOpR15 = {128'(resizzeR9[99:0]), binOpR14[255:128] * binOpR14[127:0]};
  assign resizzeR13 = binOpR15[255:128] >> binOpR15[127:0];
  assign res = (gzdLLziMainzidev6[0] == 1'h1) ? resizzeR13[0] : resizzeR8[0];
endmodule

module zdLLziMainzidev11 (input logic [99:0] arg0,
  input logic [6:0] arg1,
  output logic [0:0] res);
  logic [6:0] resizze;
  logic [255:0] binOp;
  logic [6:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [107:0] gzdLLziMainzidev10;
  logic [99:0] gMainzix2;
  logic [99:0] callRes;
  logic [99:0] resizzeR2;
  logic [6:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [6:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR6;
  logic [6:0] resizzeR7;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [127:0] resizzeR8;
  logic [6:0] resizzeR9;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [127:0] resizzeR10;
  logic [107:0] gzdLLziMainzidev9;
  logic [99:0] resizzeR11;
  logic [6:0] resizzeR12;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [127:0] resizzeR13;
  logic [6:0] resizzeR14;
  logic [255:0] binOpR14;
  logic [255:0] binOpR15;
  logic [127:0] resizzeR15;
  logic [6:0] resizzeR16;
  logic [255:0] binOpR16;
  logic [255:0] binOpR17;
  logic [255:0] binOpR18;
  logic [255:0] binOpR19;
  logic [127:0] resizzeR17;
  assign resizze = arg1;
  assign binOp = {128'(resizze[6:0]), 128'h00000000000000000000000000000031};
  assign resizzeR1 = arg1;
  assign binOpR1 = {128'(resizzeR1[6:0]), 128'h00000000000000000000000000000031};
  assign gzdLLziMainzidev10 = {arg0, arg1, binOpR1[255:128] < binOpR1[127:0]};
  assign gMainzix2 = gzdLLziMainzidev10[107:8];
  Mainzix2  Mainzix2 (gMainzix2[99:0], callRes);
  assign resizzeR2 = callRes;
  assign resizzeR3 = gzdLLziMainzidev10[7:1];
  assign binOpR2 = {128'(resizzeR3[6:0]), 128'h00000000000000000000000000000031};
  assign binOpR3 = {binOpR2[255:128] - binOpR2[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[6:0];
  assign binOpR4 = {128'(resizzeR5[6:0]), 128'h00000000000000000000000000000002};
  assign binOpR5 = {binOpR4[255:128] * binOpR4[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR6 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR7 = resizzeR6[6:0];
  assign binOpR6 = {128'(resizzeR7[6:0]), 128'h00000000000000000000000000000001};
  assign binOpR7 = {binOpR6[255:128] + binOpR6[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR8 = binOpR7[255:128] % binOpR7[127:0];
  assign resizzeR9 = resizzeR8[6:0];
  assign binOpR8 = {128'h00000000000000000000000000000064, 128'(resizzeR9[6:0])};
  assign binOpR9 = {binOpR8[255:128] - binOpR8[127:0], 128'h00000000000000000000000000000001};
  assign binOpR10 = {binOpR9[255:128] - binOpR9[127:0], 128'h00000000000000000000000000000001};
  assign binOpR11 = {128'(resizzeR2[99:0]), binOpR10[255:128] * binOpR10[127:0]};
  assign resizzeR10 = binOpR11[255:128] >> binOpR11[127:0];
  assign gzdLLziMainzidev9 = {arg0, arg1, binOp[255:128] < binOp[127:0]};
  assign resizzeR11 = gzdLLziMainzidev9[107:8];
  assign resizzeR12 = gzdLLziMainzidev9[7:1];
  assign binOpR12 = {128'(resizzeR12[6:0]), 128'h00000000000000000000000000000002};
  assign binOpR13 = {binOpR12[255:128] * binOpR12[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR13 = binOpR13[255:128] % binOpR13[127:0];
  assign resizzeR14 = resizzeR13[6:0];
  assign binOpR14 = {128'(resizzeR14[6:0]), 128'h00000000000000000000000000000001};
  assign binOpR15 = {binOpR14[255:128] + binOpR14[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR15 = binOpR15[255:128] % binOpR15[127:0];
  assign resizzeR16 = resizzeR15[6:0];
  assign binOpR16 = {128'h00000000000000000000000000000064, 128'(resizzeR16[6:0])};
  assign binOpR17 = {binOpR16[255:128] - binOpR16[127:0], 128'h00000000000000000000000000000001};
  assign binOpR18 = {binOpR17[255:128] - binOpR17[127:0], 128'h00000000000000000000000000000001};
  assign binOpR19 = {128'(resizzeR11[99:0]), binOpR18[255:128] * binOpR18[127:0]};
  assign resizzeR17 = binOpR19[255:128] >> binOpR19[127:0];
  assign res = (gzdLLziMainzidev9[0] == 1'h1) ? resizzeR17[0] : resizzeR10[0];
endmodule

module Mainzix2 (input logic [99:0] arg0,
  output logic [99:0] res);
  logic [199:0] binOp;
  assign binOp = {arg0, 100'h0000000000000000000000002};
  assign res = binOp[199:100] * binOp[99:0];
endmodule

module ReWireziPreludezinot (input logic [0:0] arg0,
  output logic [0:0] res);
  logic [0:0] lit;
  assign lit = arg0;
  assign res = (lit[0] == 1'h1) ? 1'h0 : 1'h1;
endmodule