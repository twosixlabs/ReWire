module top_level ();
  logic [0:0] __continue;
  assign __continue = 1'h1;
endmodule