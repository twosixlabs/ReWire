module top_level (input logic [63:0] __in0,
  input logic [63:0] __in1,
  output logic [63:0] __out0,
  output logic [63:0] __out1);
  logic [127:0] zll_main_loop3_in;
  logic [127:0] zll_main_compute151_in;
  logic [127:0] zll_main_compute344_in;
  logic [127:0] zll_main_compute214_in;
  logic [127:0] zll_main_compute387_in;
  logic [127:0] zll_main_compute212_in;
  logic [130:0] zll_main_compute144_in;
  logic [133:0] zll_main_compute375_in;
  logic [5:0] zll_main_compute410_in;
  logic [2:0] zll_main_compute410_out;
  logic [136:0] zll_main_compute324_in;
  logic [70:0] zll_main_compute290_in;
  logic [6:0] zll_main_compute382_in;
  logic [6:0] zll_main_compute79_in;
  logic [5:0] zll_main_compute411_in;
  logic [2:0] zll_main_compute411_out;
  logic [3:0] id_in;
  logic [133:0] zll_main_compute4_in;
  logic [136:0] zll_main_compute126_in;
  logic [7:0] zll_main_compute126_out;
  logic [136:0] zll_main_compute126_inR1;
  logic [7:0] zll_main_compute126_outR1;
  logic [136:0] zll_main_compute126_inR2;
  logic [7:0] zll_main_compute126_outR2;
  logic [136:0] zll_main_compute126_inR3;
  logic [7:0] zll_main_compute126_outR3;
  logic [136:0] zll_main_compute126_inR4;
  logic [7:0] zll_main_compute126_outR4;
  logic [136:0] zll_main_compute126_inR5;
  logic [7:0] zll_main_compute126_outR5;
  logic [136:0] zll_main_compute126_inR6;
  logic [7:0] zll_main_compute126_outR6;
  logic [136:0] zll_main_compute126_inR7;
  logic [7:0] zll_main_compute126_outR7;
  logic [127:0] zll_main_compute284_in;
  logic [127:0] zll_main_compute287_in;
  logic [127:0] zll_main_compute89_in;
  logic [130:0] zll_main_compute323_in;
  logic [130:0] zll_main_compute398_in;
  logic [133:0] zll_main_compute265_in;
  logic [5:0] zll_main_compute410_inR1;
  logic [2:0] zll_main_compute410_outR1;
  logic [136:0] zll_main_compute75_in;
  logic [70:0] zll_main_compute386_in;
  logic [2:0] zll_main_compute386_out;
  logic [136:0] zll_main_compute263_in;
  logic [139:0] zll_main_compute232_in;
  logic [7:0] zll_main_compute232_out;
  logic [139:0] zll_main_compute232_inR1;
  logic [7:0] zll_main_compute232_outR1;
  logic [139:0] zll_main_compute232_inR2;
  logic [7:0] zll_main_compute232_outR2;
  logic [139:0] zll_main_compute232_inR3;
  logic [7:0] zll_main_compute232_outR3;
  logic [139:0] zll_main_compute232_inR4;
  logic [7:0] zll_main_compute232_outR4;
  logic [139:0] zll_main_compute232_inR5;
  logic [7:0] zll_main_compute232_outR5;
  logic [139:0] zll_main_compute232_inR6;
  logic [7:0] zll_main_compute232_outR6;
  logic [139:0] zll_main_compute232_inR7;
  logic [7:0] zll_main_compute232_outR7;
  logic [127:0] zll_main_compute132_in;
  logic [127:0] zll_main_compute417_in;
  logic [127:0] zll_main_compute330_in;
  logic [127:0] zll_main_compute42_in;
  logic [127:0] zll_main_compute403_in;
  logic [127:0] zll_main_compute229_in;
  logic [130:0] zll_main_compute73_in;
  logic [130:0] zll_main_compute58_in;
  logic [133:0] zll_main_compute159_in;
  logic [5:0] zll_main_compute410_inR2;
  logic [2:0] zll_main_compute410_outR2;
  logic [136:0] zll_main_compute420_in;
  logic [70:0] zll_main_compute386_inR1;
  logic [2:0] zll_main_compute386_outR1;
  logic [133:0] zll_main_compute181_in;
  logic [136:0] zll_main_compute41_in;
  logic [7:0] zll_main_compute41_out;
  logic [136:0] zll_main_compute41_inR1;
  logic [7:0] zll_main_compute41_outR1;
  logic [136:0] zll_main_compute41_inR2;
  logic [7:0] zll_main_compute41_outR2;
  logic [136:0] zll_main_compute41_inR3;
  logic [7:0] zll_main_compute41_outR3;
  logic [136:0] zll_main_compute41_inR4;
  logic [7:0] zll_main_compute41_outR4;
  logic [136:0] zll_main_compute41_inR5;
  logic [7:0] zll_main_compute41_outR5;
  logic [136:0] zll_main_compute41_inR6;
  logic [7:0] zll_main_compute41_outR6;
  logic [136:0] zll_main_compute41_inR7;
  logic [7:0] zll_main_compute41_outR7;
  logic [127:0] zll_main_compute277_in;
  logic [127:0] zll_main_compute111_in;
  logic [127:0] zll_main_compute32_in;
  logic [130:0] zll_main_compute405_in;
  logic [130:0] zll_main_compute367_in;
  logic [133:0] zll_main_compute43_in;
  logic [5:0] zll_main_compute410_inR3;
  logic [2:0] zll_main_compute410_outR3;
  logic [136:0] zll_main_compute427_in;
  logic [70:0] zll_main_compute386_inR2;
  logic [2:0] zll_main_compute386_outR2;
  logic [136:0] zll_main_compute447_in;
  logic [139:0] zll_main_compute215_in;
  logic [7:0] zll_main_compute215_out;
  logic [139:0] zll_main_compute215_inR1;
  logic [7:0] zll_main_compute215_outR1;
  logic [139:0] zll_main_compute215_inR2;
  logic [7:0] zll_main_compute215_outR2;
  logic [139:0] zll_main_compute215_inR3;
  logic [7:0] zll_main_compute215_outR3;
  logic [139:0] zll_main_compute215_inR4;
  logic [7:0] zll_main_compute215_outR4;
  logic [139:0] zll_main_compute215_inR5;
  logic [7:0] zll_main_compute215_outR5;
  logic [139:0] zll_main_compute215_inR6;
  logic [7:0] zll_main_compute215_outR6;
  logic [139:0] zll_main_compute215_inR7;
  logic [7:0] zll_main_compute215_outR7;
  logic [127:0] zll_main_compute154_in;
  logic [127:0] zll_main_compute117_in;
  logic [127:0] zll_main_compute329_in;
  logic [127:0] zll_main_compute205_in;
  logic [127:0] zll_main_compute278_in;
  logic [130:0] zll_main_compute195_in;
  logic [130:0] zll_main_compute254_in;
  logic [133:0] zll_main_compute90_in;
  logic [136:0] zll_main_compute238_in;
  logic [7:0] zll_main_compute238_out;
  logic [136:0] zll_main_compute238_inR1;
  logic [7:0] zll_main_compute238_outR1;
  logic [136:0] zll_main_compute238_inR2;
  logic [7:0] zll_main_compute238_outR2;
  logic [136:0] zll_main_compute238_inR3;
  logic [7:0] zll_main_compute238_outR3;
  logic [136:0] zll_main_compute238_inR4;
  logic [7:0] zll_main_compute238_outR4;
  logic [136:0] zll_main_compute238_inR5;
  logic [7:0] zll_main_compute238_outR5;
  logic [136:0] zll_main_compute238_inR6;
  logic [7:0] zll_main_compute238_outR6;
  logic [136:0] zll_main_compute238_inR7;
  logic [7:0] zll_main_compute238_outR7;
  logic [127:0] zll_main_compute209_in;
  logic [127:0] zll_main_compute28_in;
  logic [127:0] zll_main_compute436_in;
  logic [130:0] zll_main_compute280_in;
  logic [133:0] zll_main_compute82_in;
  logic [5:0] zll_main_compute410_inR4;
  logic [2:0] zll_main_compute410_outR4;
  logic [136:0] zll_main_compute452_in;
  logic [70:0] zll_main_compute173_in;
  logic [6:0] zll_main_compute270_in;
  logic [2:0] zll_main_compute270_out;
  logic [3:0] id_inR1;
  logic [136:0] zll_main_compute39_in;
  logic [139:0] zll_main_compute187_in;
  logic [7:0] zll_main_compute187_out;
  logic [139:0] zll_main_compute187_inR1;
  logic [7:0] zll_main_compute187_outR1;
  logic [139:0] zll_main_compute187_inR2;
  logic [7:0] zll_main_compute187_outR2;
  logic [139:0] zll_main_compute187_inR3;
  logic [7:0] zll_main_compute187_outR3;
  logic [139:0] zll_main_compute187_inR4;
  logic [7:0] zll_main_compute187_outR4;
  logic [139:0] zll_main_compute187_inR5;
  logic [7:0] zll_main_compute187_outR5;
  logic [139:0] zll_main_compute187_inR6;
  logic [7:0] zll_main_compute187_outR6;
  logic [139:0] zll_main_compute187_inR7;
  logic [7:0] zll_main_compute187_outR7;
  logic [127:0] zll_main_compute258_in;
  logic [127:0] id_inR2;
  logic [128:0] zll_main_loop2_in;
  logic [128:0] zll_main_loop_in;
  logic [0:0] __padding;
  assign zll_main_loop3_in = {__in0, __in1};
  assign zll_main_compute151_in = zll_main_loop3_in[127:0];
  assign zll_main_compute344_in = zll_main_compute151_in[127:0];
  assign zll_main_compute214_in = {zll_main_compute344_in[127:64], zll_main_compute344_in[63:0]};
  assign zll_main_compute387_in = {zll_main_compute214_in[127:64], zll_main_compute214_in[63:0]};
  assign zll_main_compute212_in = zll_main_compute387_in[127:0];
  assign zll_main_compute144_in = {zll_main_compute212_in[127:64], zll_main_compute212_in[63:0], 3'h1};
  assign zll_main_compute375_in = {zll_main_compute144_in[130:67], zll_main_compute144_in[66:3], zll_main_compute144_in[2:0], 3'h2};
  assign zll_main_compute410_in = {3'h7, zll_main_compute375_in[2:0]};
  ZLL_Main_compute410  inst (zll_main_compute410_in[5:3], zll_main_compute410_in[2:0], zll_main_compute410_out);
  assign zll_main_compute324_in = {zll_main_compute375_in[2:0], zll_main_compute375_in[133:70], zll_main_compute375_in[69:6], zll_main_compute375_in[5:3], zll_main_compute410_out};
  assign zll_main_compute290_in = {zll_main_compute324_in[2:0], zll_main_compute324_in[133:70], zll_main_compute324_in[5:3], 1'h0};
  assign zll_main_compute382_in = {zll_main_compute290_in[70:68], zll_main_compute290_in[3:1], 1'h0};
  assign zll_main_compute79_in = {zll_main_compute382_in[6:4], zll_main_compute382_in[3:1], zll_main_compute382_in[0]};
  assign zll_main_compute411_in = {zll_main_compute79_in[6:4], zll_main_compute79_in[3:1]};
  ZLL_Main_compute411  instR1 (zll_main_compute411_in[5:3], zll_main_compute411_in[2:0], zll_main_compute411_out);
  assign id_in = {zll_main_compute290_in[70:68], zll_main_compute290_in[0]};
  assign zll_main_compute4_in = {zll_main_compute324_in[136:134], zll_main_compute324_in[133:70], zll_main_compute324_in[69:6], (id_in[0] == 1'h1) ? id_in[3:1] : zll_main_compute411_out};
  assign zll_main_compute126_in = {zll_main_compute4_in[133:131], zll_main_compute4_in[130:67], zll_main_compute4_in[2:0], zll_main_compute4_in[66:3], 3'h0};
  ZLL_Main_compute126  instR2 (zll_main_compute126_in[136:134], zll_main_compute126_in[133:70], zll_main_compute126_in[69:67], zll_main_compute126_in[66:3], zll_main_compute126_in[2:0], zll_main_compute126_out);
  assign zll_main_compute126_inR1 = {zll_main_compute4_in[133:131], zll_main_compute4_in[130:67], zll_main_compute4_in[2:0], zll_main_compute4_in[66:3], 3'h1};
  ZLL_Main_compute126  instR3 (zll_main_compute126_inR1[136:134], zll_main_compute126_inR1[133:70], zll_main_compute126_inR1[69:67], zll_main_compute126_inR1[66:3], zll_main_compute126_inR1[2:0], zll_main_compute126_outR1);
  assign zll_main_compute126_inR2 = {zll_main_compute4_in[133:131], zll_main_compute4_in[130:67], zll_main_compute4_in[2:0], zll_main_compute4_in[66:3], 3'h2};
  ZLL_Main_compute126  instR4 (zll_main_compute126_inR2[136:134], zll_main_compute126_inR2[133:70], zll_main_compute126_inR2[69:67], zll_main_compute126_inR2[66:3], zll_main_compute126_inR2[2:0], zll_main_compute126_outR2);
  assign zll_main_compute126_inR3 = {zll_main_compute4_in[133:131], zll_main_compute4_in[130:67], zll_main_compute4_in[2:0], zll_main_compute4_in[66:3], 3'h3};
  ZLL_Main_compute126  instR5 (zll_main_compute126_inR3[136:134], zll_main_compute126_inR3[133:70], zll_main_compute126_inR3[69:67], zll_main_compute126_inR3[66:3], zll_main_compute126_inR3[2:0], zll_main_compute126_outR3);
  assign zll_main_compute126_inR4 = {zll_main_compute4_in[133:131], zll_main_compute4_in[130:67], zll_main_compute4_in[2:0], zll_main_compute4_in[66:3], 3'h4};
  ZLL_Main_compute126  instR6 (zll_main_compute126_inR4[136:134], zll_main_compute126_inR4[133:70], zll_main_compute126_inR4[69:67], zll_main_compute126_inR4[66:3], zll_main_compute126_inR4[2:0], zll_main_compute126_outR4);
  assign zll_main_compute126_inR5 = {zll_main_compute4_in[133:131], zll_main_compute4_in[130:67], zll_main_compute4_in[2:0], zll_main_compute4_in[66:3], 3'h5};
  ZLL_Main_compute126  instR7 (zll_main_compute126_inR5[136:134], zll_main_compute126_inR5[133:70], zll_main_compute126_inR5[69:67], zll_main_compute126_inR5[66:3], zll_main_compute126_inR5[2:0], zll_main_compute126_outR5);
  assign zll_main_compute126_inR6 = {zll_main_compute4_in[133:131], zll_main_compute4_in[130:67], zll_main_compute4_in[2:0], zll_main_compute4_in[66:3], 3'h6};
  ZLL_Main_compute126  instR8 (zll_main_compute126_inR6[136:134], zll_main_compute126_inR6[133:70], zll_main_compute126_inR6[69:67], zll_main_compute126_inR6[66:3], zll_main_compute126_inR6[2:0], zll_main_compute126_outR6);
  assign zll_main_compute126_inR7 = {zll_main_compute4_in[133:131], zll_main_compute4_in[130:67], zll_main_compute4_in[2:0], zll_main_compute4_in[66:3], 3'h7};
  ZLL_Main_compute126  instR9 (zll_main_compute126_inR7[136:134], zll_main_compute126_inR7[133:70], zll_main_compute126_inR7[69:67], zll_main_compute126_inR7[66:3], zll_main_compute126_inR7[2:0], zll_main_compute126_outR7);
  assign zll_main_compute284_in = {zll_main_compute344_in[127:64], zll_main_compute344_in[63:0]};
  assign zll_main_compute287_in = {zll_main_compute284_in[127:64], zll_main_compute284_in[63:0]};
  assign zll_main_compute89_in = zll_main_compute287_in[127:0];
  assign zll_main_compute323_in = {zll_main_compute89_in[127:64], zll_main_compute89_in[63:0], 3'h1};
  assign zll_main_compute398_in = {zll_main_compute323_in[2:0], zll_main_compute323_in[130:67], zll_main_compute323_in[66:3]};
  assign zll_main_compute265_in = {zll_main_compute398_in[130:128], zll_main_compute398_in[127:64], zll_main_compute398_in[63:0], 3'h2};
  assign zll_main_compute410_inR1 = {3'h7, zll_main_compute265_in[2:0]};
  ZLL_Main_compute410  instR10 (zll_main_compute410_inR1[5:3], zll_main_compute410_inR1[2:0], zll_main_compute410_outR1);
  assign zll_main_compute75_in = {zll_main_compute265_in[133:131], zll_main_compute265_in[2:0], zll_main_compute265_in[130:67], zll_main_compute265_in[66:3], zll_main_compute410_outR1};
  assign zll_main_compute386_in = {zll_main_compute75_in[136:134], zll_main_compute75_in[2:0], zll_main_compute75_in[130:67], 1'h0};
  ZLL_Main_compute386  instR11 (zll_main_compute386_in[70:68], zll_main_compute386_in[67:65], zll_main_compute386_in[64:1], zll_main_compute386_in[0], zll_main_compute386_out);
  assign zll_main_compute263_in = {zll_main_compute75_in[136:134], zll_main_compute75_in[133:131], zll_main_compute75_in[130:67], zll_main_compute75_in[66:3], zll_main_compute386_out};
  assign zll_main_compute232_in = {zll_main_compute263_in[136:134], zll_main_compute263_in[133:131], zll_main_compute263_in[130:67], zll_main_compute263_in[2:0], zll_main_compute263_in[66:3], 3'h0};
  ZLL_Main_compute232  instR12 (zll_main_compute232_in[139:137], zll_main_compute232_in[136:134], zll_main_compute232_in[133:70], zll_main_compute232_in[69:67], zll_main_compute232_in[66:3], zll_main_compute232_in[2:0], zll_main_compute232_out);
  assign zll_main_compute232_inR1 = {zll_main_compute263_in[136:134], zll_main_compute263_in[133:131], zll_main_compute263_in[130:67], zll_main_compute263_in[2:0], zll_main_compute263_in[66:3], 3'h1};
  ZLL_Main_compute232  instR13 (zll_main_compute232_inR1[139:137], zll_main_compute232_inR1[136:134], zll_main_compute232_inR1[133:70], zll_main_compute232_inR1[69:67], zll_main_compute232_inR1[66:3], zll_main_compute232_inR1[2:0], zll_main_compute232_outR1);
  assign zll_main_compute232_inR2 = {zll_main_compute263_in[136:134], zll_main_compute263_in[133:131], zll_main_compute263_in[130:67], zll_main_compute263_in[2:0], zll_main_compute263_in[66:3], 3'h2};
  ZLL_Main_compute232  instR14 (zll_main_compute232_inR2[139:137], zll_main_compute232_inR2[136:134], zll_main_compute232_inR2[133:70], zll_main_compute232_inR2[69:67], zll_main_compute232_inR2[66:3], zll_main_compute232_inR2[2:0], zll_main_compute232_outR2);
  assign zll_main_compute232_inR3 = {zll_main_compute263_in[136:134], zll_main_compute263_in[133:131], zll_main_compute263_in[130:67], zll_main_compute263_in[2:0], zll_main_compute263_in[66:3], 3'h3};
  ZLL_Main_compute232  instR15 (zll_main_compute232_inR3[139:137], zll_main_compute232_inR3[136:134], zll_main_compute232_inR3[133:70], zll_main_compute232_inR3[69:67], zll_main_compute232_inR3[66:3], zll_main_compute232_inR3[2:0], zll_main_compute232_outR3);
  assign zll_main_compute232_inR4 = {zll_main_compute263_in[136:134], zll_main_compute263_in[133:131], zll_main_compute263_in[130:67], zll_main_compute263_in[2:0], zll_main_compute263_in[66:3], 3'h4};
  ZLL_Main_compute232  instR16 (zll_main_compute232_inR4[139:137], zll_main_compute232_inR4[136:134], zll_main_compute232_inR4[133:70], zll_main_compute232_inR4[69:67], zll_main_compute232_inR4[66:3], zll_main_compute232_inR4[2:0], zll_main_compute232_outR4);
  assign zll_main_compute232_inR5 = {zll_main_compute263_in[136:134], zll_main_compute263_in[133:131], zll_main_compute263_in[130:67], zll_main_compute263_in[2:0], zll_main_compute263_in[66:3], 3'h5};
  ZLL_Main_compute232  instR17 (zll_main_compute232_inR5[139:137], zll_main_compute232_inR5[136:134], zll_main_compute232_inR5[133:70], zll_main_compute232_inR5[69:67], zll_main_compute232_inR5[66:3], zll_main_compute232_inR5[2:0], zll_main_compute232_outR5);
  assign zll_main_compute232_inR6 = {zll_main_compute263_in[136:134], zll_main_compute263_in[133:131], zll_main_compute263_in[130:67], zll_main_compute263_in[2:0], zll_main_compute263_in[66:3], 3'h6};
  ZLL_Main_compute232  instR18 (zll_main_compute232_inR6[139:137], zll_main_compute232_inR6[136:134], zll_main_compute232_inR6[133:70], zll_main_compute232_inR6[69:67], zll_main_compute232_inR6[66:3], zll_main_compute232_inR6[2:0], zll_main_compute232_outR6);
  assign zll_main_compute232_inR7 = {zll_main_compute263_in[136:134], zll_main_compute263_in[133:131], zll_main_compute263_in[130:67], zll_main_compute263_in[2:0], zll_main_compute263_in[66:3], 3'h7};
  ZLL_Main_compute232  instR19 (zll_main_compute232_inR7[139:137], zll_main_compute232_inR7[136:134], zll_main_compute232_inR7[133:70], zll_main_compute232_inR7[69:67], zll_main_compute232_inR7[66:3], zll_main_compute232_inR7[2:0], zll_main_compute232_outR7);
  assign zll_main_compute132_in = {{zll_main_compute126_out, zll_main_compute126_outR1, zll_main_compute126_outR2, zll_main_compute126_outR3, zll_main_compute126_outR4, zll_main_compute126_outR5, zll_main_compute126_outR6, zll_main_compute126_outR7}, {zll_main_compute232_out, zll_main_compute232_outR1, zll_main_compute232_outR2, zll_main_compute232_outR3, zll_main_compute232_outR4, zll_main_compute232_outR5, zll_main_compute232_outR6, zll_main_compute232_outR7}};
  assign zll_main_compute417_in = zll_main_compute132_in[127:0];
  assign zll_main_compute330_in = {zll_main_compute417_in[63:0], zll_main_compute417_in[127:64]};
  assign zll_main_compute42_in = {zll_main_compute330_in[127:64], zll_main_compute330_in[63:0]};
  assign zll_main_compute403_in = zll_main_compute42_in[127:0];
  assign zll_main_compute229_in = {zll_main_compute403_in[63:0], zll_main_compute403_in[127:64]};
  assign zll_main_compute73_in = {zll_main_compute229_in[127:64], zll_main_compute229_in[63:0], 3'h1};
  assign zll_main_compute58_in = {zll_main_compute73_in[130:67], zll_main_compute73_in[2:0], zll_main_compute73_in[66:3]};
  assign zll_main_compute159_in = {zll_main_compute58_in[130:67], zll_main_compute58_in[66:64], zll_main_compute58_in[63:0], 3'h2};
  assign zll_main_compute410_inR2 = {3'h7, zll_main_compute159_in[2:0]};
  ZLL_Main_compute410  instR20 (zll_main_compute410_inR2[5:3], zll_main_compute410_inR2[2:0], zll_main_compute410_outR2);
  assign zll_main_compute420_in = {zll_main_compute159_in[2:0], zll_main_compute159_in[133:70], zll_main_compute159_in[69:67], zll_main_compute159_in[66:3], zll_main_compute410_outR2};
  assign zll_main_compute386_inR1 = {zll_main_compute420_in[69:67], zll_main_compute420_in[2:0], zll_main_compute420_in[66:3], 1'h0};
  ZLL_Main_compute386  instR21 (zll_main_compute386_inR1[70:68], zll_main_compute386_inR1[67:65], zll_main_compute386_inR1[64:1], zll_main_compute386_inR1[0], zll_main_compute386_outR1);
  assign zll_main_compute181_in = {zll_main_compute420_in[136:134], zll_main_compute420_in[133:70], zll_main_compute420_in[66:3], zll_main_compute386_outR1};
  assign zll_main_compute41_in = {zll_main_compute181_in[133:131], zll_main_compute181_in[130:67], zll_main_compute181_in[2:0], zll_main_compute181_in[66:3], 3'h0};
  ZLL_Main_compute41  instR22 (zll_main_compute41_in[136:134], zll_main_compute41_in[133:70], zll_main_compute41_in[69:67], zll_main_compute41_in[66:3], zll_main_compute41_in[2:0], zll_main_compute41_out);
  assign zll_main_compute41_inR1 = {zll_main_compute181_in[133:131], zll_main_compute181_in[130:67], zll_main_compute181_in[2:0], zll_main_compute181_in[66:3], 3'h1};
  ZLL_Main_compute41  instR23 (zll_main_compute41_inR1[136:134], zll_main_compute41_inR1[133:70], zll_main_compute41_inR1[69:67], zll_main_compute41_inR1[66:3], zll_main_compute41_inR1[2:0], zll_main_compute41_outR1);
  assign zll_main_compute41_inR2 = {zll_main_compute181_in[133:131], zll_main_compute181_in[130:67], zll_main_compute181_in[2:0], zll_main_compute181_in[66:3], 3'h2};
  ZLL_Main_compute41  instR24 (zll_main_compute41_inR2[136:134], zll_main_compute41_inR2[133:70], zll_main_compute41_inR2[69:67], zll_main_compute41_inR2[66:3], zll_main_compute41_inR2[2:0], zll_main_compute41_outR2);
  assign zll_main_compute41_inR3 = {zll_main_compute181_in[133:131], zll_main_compute181_in[130:67], zll_main_compute181_in[2:0], zll_main_compute181_in[66:3], 3'h3};
  ZLL_Main_compute41  instR25 (zll_main_compute41_inR3[136:134], zll_main_compute41_inR3[133:70], zll_main_compute41_inR3[69:67], zll_main_compute41_inR3[66:3], zll_main_compute41_inR3[2:0], zll_main_compute41_outR3);
  assign zll_main_compute41_inR4 = {zll_main_compute181_in[133:131], zll_main_compute181_in[130:67], zll_main_compute181_in[2:0], zll_main_compute181_in[66:3], 3'h4};
  ZLL_Main_compute41  instR26 (zll_main_compute41_inR4[136:134], zll_main_compute41_inR4[133:70], zll_main_compute41_inR4[69:67], zll_main_compute41_inR4[66:3], zll_main_compute41_inR4[2:0], zll_main_compute41_outR4);
  assign zll_main_compute41_inR5 = {zll_main_compute181_in[133:131], zll_main_compute181_in[130:67], zll_main_compute181_in[2:0], zll_main_compute181_in[66:3], 3'h5};
  ZLL_Main_compute41  instR27 (zll_main_compute41_inR5[136:134], zll_main_compute41_inR5[133:70], zll_main_compute41_inR5[69:67], zll_main_compute41_inR5[66:3], zll_main_compute41_inR5[2:0], zll_main_compute41_outR5);
  assign zll_main_compute41_inR6 = {zll_main_compute181_in[133:131], zll_main_compute181_in[130:67], zll_main_compute181_in[2:0], zll_main_compute181_in[66:3], 3'h6};
  ZLL_Main_compute41  instR28 (zll_main_compute41_inR6[136:134], zll_main_compute41_inR6[133:70], zll_main_compute41_inR6[69:67], zll_main_compute41_inR6[66:3], zll_main_compute41_inR6[2:0], zll_main_compute41_outR6);
  assign zll_main_compute41_inR7 = {zll_main_compute181_in[133:131], zll_main_compute181_in[130:67], zll_main_compute181_in[2:0], zll_main_compute181_in[66:3], 3'h7};
  ZLL_Main_compute41  instR29 (zll_main_compute41_inR7[136:134], zll_main_compute41_inR7[133:70], zll_main_compute41_inR7[69:67], zll_main_compute41_inR7[66:3], zll_main_compute41_inR7[2:0], zll_main_compute41_outR7);
  assign zll_main_compute277_in = {zll_main_compute417_in[63:0], zll_main_compute417_in[127:64]};
  assign zll_main_compute111_in = {zll_main_compute277_in[127:64], zll_main_compute277_in[63:0]};
  assign zll_main_compute32_in = zll_main_compute111_in[127:0];
  assign zll_main_compute405_in = {zll_main_compute32_in[127:64], zll_main_compute32_in[63:0], 3'h1};
  assign zll_main_compute367_in = {zll_main_compute405_in[2:0], zll_main_compute405_in[130:67], zll_main_compute405_in[66:3]};
  assign zll_main_compute43_in = {zll_main_compute367_in[130:128], zll_main_compute367_in[127:64], zll_main_compute367_in[63:0], 3'h2};
  assign zll_main_compute410_inR3 = {3'h7, zll_main_compute43_in[2:0]};
  ZLL_Main_compute410  instR30 (zll_main_compute410_inR3[5:3], zll_main_compute410_inR3[2:0], zll_main_compute410_outR3);
  assign zll_main_compute427_in = {zll_main_compute43_in[2:0], zll_main_compute43_in[133:131], zll_main_compute43_in[130:67], zll_main_compute43_in[66:3], zll_main_compute410_outR3};
  assign zll_main_compute386_inR2 = {zll_main_compute427_in[133:131], zll_main_compute427_in[2:0], zll_main_compute427_in[130:67], 1'h0};
  ZLL_Main_compute386  instR31 (zll_main_compute386_inR2[70:68], zll_main_compute386_inR2[67:65], zll_main_compute386_inR2[64:1], zll_main_compute386_inR2[0], zll_main_compute386_outR2);
  assign zll_main_compute447_in = {zll_main_compute427_in[136:134], zll_main_compute427_in[133:131], zll_main_compute427_in[130:67], zll_main_compute427_in[66:3], zll_main_compute386_outR2};
  assign zll_main_compute215_in = {zll_main_compute447_in[136:134], zll_main_compute447_in[133:131], zll_main_compute447_in[130:67], zll_main_compute447_in[66:3], zll_main_compute447_in[2:0], 3'h0};
  ZLL_Main_compute215  instR32 (zll_main_compute215_in[139:137], zll_main_compute215_in[136:134], zll_main_compute215_in[133:70], zll_main_compute215_in[69:6], zll_main_compute215_in[5:3], zll_main_compute215_in[2:0], zll_main_compute215_out);
  assign zll_main_compute215_inR1 = {zll_main_compute447_in[136:134], zll_main_compute447_in[133:131], zll_main_compute447_in[130:67], zll_main_compute447_in[66:3], zll_main_compute447_in[2:0], 3'h1};
  ZLL_Main_compute215  instR33 (zll_main_compute215_inR1[139:137], zll_main_compute215_inR1[136:134], zll_main_compute215_inR1[133:70], zll_main_compute215_inR1[69:6], zll_main_compute215_inR1[5:3], zll_main_compute215_inR1[2:0], zll_main_compute215_outR1);
  assign zll_main_compute215_inR2 = {zll_main_compute447_in[136:134], zll_main_compute447_in[133:131], zll_main_compute447_in[130:67], zll_main_compute447_in[66:3], zll_main_compute447_in[2:0], 3'h2};
  ZLL_Main_compute215  instR34 (zll_main_compute215_inR2[139:137], zll_main_compute215_inR2[136:134], zll_main_compute215_inR2[133:70], zll_main_compute215_inR2[69:6], zll_main_compute215_inR2[5:3], zll_main_compute215_inR2[2:0], zll_main_compute215_outR2);
  assign zll_main_compute215_inR3 = {zll_main_compute447_in[136:134], zll_main_compute447_in[133:131], zll_main_compute447_in[130:67], zll_main_compute447_in[66:3], zll_main_compute447_in[2:0], 3'h3};
  ZLL_Main_compute215  instR35 (zll_main_compute215_inR3[139:137], zll_main_compute215_inR3[136:134], zll_main_compute215_inR3[133:70], zll_main_compute215_inR3[69:6], zll_main_compute215_inR3[5:3], zll_main_compute215_inR3[2:0], zll_main_compute215_outR3);
  assign zll_main_compute215_inR4 = {zll_main_compute447_in[136:134], zll_main_compute447_in[133:131], zll_main_compute447_in[130:67], zll_main_compute447_in[66:3], zll_main_compute447_in[2:0], 3'h4};
  ZLL_Main_compute215  instR36 (zll_main_compute215_inR4[139:137], zll_main_compute215_inR4[136:134], zll_main_compute215_inR4[133:70], zll_main_compute215_inR4[69:6], zll_main_compute215_inR4[5:3], zll_main_compute215_inR4[2:0], zll_main_compute215_outR4);
  assign zll_main_compute215_inR5 = {zll_main_compute447_in[136:134], zll_main_compute447_in[133:131], zll_main_compute447_in[130:67], zll_main_compute447_in[66:3], zll_main_compute447_in[2:0], 3'h5};
  ZLL_Main_compute215  instR37 (zll_main_compute215_inR5[139:137], zll_main_compute215_inR5[136:134], zll_main_compute215_inR5[133:70], zll_main_compute215_inR5[69:6], zll_main_compute215_inR5[5:3], zll_main_compute215_inR5[2:0], zll_main_compute215_outR5);
  assign zll_main_compute215_inR6 = {zll_main_compute447_in[136:134], zll_main_compute447_in[133:131], zll_main_compute447_in[130:67], zll_main_compute447_in[66:3], zll_main_compute447_in[2:0], 3'h6};
  ZLL_Main_compute215  instR38 (zll_main_compute215_inR6[139:137], zll_main_compute215_inR6[136:134], zll_main_compute215_inR6[133:70], zll_main_compute215_inR6[69:6], zll_main_compute215_inR6[5:3], zll_main_compute215_inR6[2:0], zll_main_compute215_outR6);
  assign zll_main_compute215_inR7 = {zll_main_compute447_in[136:134], zll_main_compute447_in[133:131], zll_main_compute447_in[130:67], zll_main_compute447_in[66:3], zll_main_compute447_in[2:0], 3'h7};
  ZLL_Main_compute215  instR39 (zll_main_compute215_inR7[139:137], zll_main_compute215_inR7[136:134], zll_main_compute215_inR7[133:70], zll_main_compute215_inR7[69:6], zll_main_compute215_inR7[5:3], zll_main_compute215_inR7[2:0], zll_main_compute215_outR7);
  assign zll_main_compute154_in = {{zll_main_compute41_out, zll_main_compute41_outR1, zll_main_compute41_outR2, zll_main_compute41_outR3, zll_main_compute41_outR4, zll_main_compute41_outR5, zll_main_compute41_outR6, zll_main_compute41_outR7}, {zll_main_compute215_out, zll_main_compute215_outR1, zll_main_compute215_outR2, zll_main_compute215_outR3, zll_main_compute215_outR4, zll_main_compute215_outR5, zll_main_compute215_outR6, zll_main_compute215_outR7}};
  assign zll_main_compute117_in = zll_main_compute154_in[127:0];
  assign zll_main_compute329_in = {zll_main_compute117_in[127:64], zll_main_compute117_in[63:0]};
  assign zll_main_compute205_in = {zll_main_compute329_in[127:64], zll_main_compute329_in[63:0]};
  assign zll_main_compute278_in = zll_main_compute205_in[127:0];
  assign zll_main_compute195_in = {zll_main_compute278_in[127:64], zll_main_compute278_in[63:0], 3'h1};
  assign zll_main_compute254_in = {zll_main_compute195_in[130:67], zll_main_compute195_in[2:0], zll_main_compute195_in[66:3]};
  assign zll_main_compute90_in = {zll_main_compute254_in[130:67], zll_main_compute254_in[66:64], zll_main_compute254_in[63:0], 3'h2};
  assign zll_main_compute238_in = {zll_main_compute90_in[133:70], zll_main_compute90_in[2:0], zll_main_compute90_in[69:67], zll_main_compute90_in[66:3], 3'h0};
  ZLL_Main_compute238  instR40 (zll_main_compute238_in[136:73], zll_main_compute238_in[72:70], zll_main_compute238_in[69:67], zll_main_compute238_in[66:3], zll_main_compute238_in[2:0], zll_main_compute238_out);
  assign zll_main_compute238_inR1 = {zll_main_compute90_in[133:70], zll_main_compute90_in[2:0], zll_main_compute90_in[69:67], zll_main_compute90_in[66:3], 3'h1};
  ZLL_Main_compute238  instR41 (zll_main_compute238_inR1[136:73], zll_main_compute238_inR1[72:70], zll_main_compute238_inR1[69:67], zll_main_compute238_inR1[66:3], zll_main_compute238_inR1[2:0], zll_main_compute238_outR1);
  assign zll_main_compute238_inR2 = {zll_main_compute90_in[133:70], zll_main_compute90_in[2:0], zll_main_compute90_in[69:67], zll_main_compute90_in[66:3], 3'h2};
  ZLL_Main_compute238  instR42 (zll_main_compute238_inR2[136:73], zll_main_compute238_inR2[72:70], zll_main_compute238_inR2[69:67], zll_main_compute238_inR2[66:3], zll_main_compute238_inR2[2:0], zll_main_compute238_outR2);
  assign zll_main_compute238_inR3 = {zll_main_compute90_in[133:70], zll_main_compute90_in[2:0], zll_main_compute90_in[69:67], zll_main_compute90_in[66:3], 3'h3};
  ZLL_Main_compute238  instR43 (zll_main_compute238_inR3[136:73], zll_main_compute238_inR3[72:70], zll_main_compute238_inR3[69:67], zll_main_compute238_inR3[66:3], zll_main_compute238_inR3[2:0], zll_main_compute238_outR3);
  assign zll_main_compute238_inR4 = {zll_main_compute90_in[133:70], zll_main_compute90_in[2:0], zll_main_compute90_in[69:67], zll_main_compute90_in[66:3], 3'h4};
  ZLL_Main_compute238  instR44 (zll_main_compute238_inR4[136:73], zll_main_compute238_inR4[72:70], zll_main_compute238_inR4[69:67], zll_main_compute238_inR4[66:3], zll_main_compute238_inR4[2:0], zll_main_compute238_outR4);
  assign zll_main_compute238_inR5 = {zll_main_compute90_in[133:70], zll_main_compute90_in[2:0], zll_main_compute90_in[69:67], zll_main_compute90_in[66:3], 3'h5};
  ZLL_Main_compute238  instR45 (zll_main_compute238_inR5[136:73], zll_main_compute238_inR5[72:70], zll_main_compute238_inR5[69:67], zll_main_compute238_inR5[66:3], zll_main_compute238_inR5[2:0], zll_main_compute238_outR5);
  assign zll_main_compute238_inR6 = {zll_main_compute90_in[133:70], zll_main_compute90_in[2:0], zll_main_compute90_in[69:67], zll_main_compute90_in[66:3], 3'h6};
  ZLL_Main_compute238  instR46 (zll_main_compute238_inR6[136:73], zll_main_compute238_inR6[72:70], zll_main_compute238_inR6[69:67], zll_main_compute238_inR6[66:3], zll_main_compute238_inR6[2:0], zll_main_compute238_outR6);
  assign zll_main_compute238_inR7 = {zll_main_compute90_in[133:70], zll_main_compute90_in[2:0], zll_main_compute90_in[69:67], zll_main_compute90_in[66:3], 3'h7};
  ZLL_Main_compute238  instR47 (zll_main_compute238_inR7[136:73], zll_main_compute238_inR7[72:70], zll_main_compute238_inR7[69:67], zll_main_compute238_inR7[66:3], zll_main_compute238_inR7[2:0], zll_main_compute238_outR7);
  assign zll_main_compute209_in = {zll_main_compute117_in[127:64], zll_main_compute117_in[63:0]};
  assign zll_main_compute28_in = {zll_main_compute209_in[127:64], zll_main_compute209_in[63:0]};
  assign zll_main_compute436_in = zll_main_compute28_in[127:0];
  assign zll_main_compute280_in = {zll_main_compute436_in[127:64], zll_main_compute436_in[63:0], 3'h1};
  assign zll_main_compute82_in = {zll_main_compute280_in[130:67], zll_main_compute280_in[66:3], zll_main_compute280_in[2:0], 3'h2};
  assign zll_main_compute410_inR4 = {3'h7, zll_main_compute82_in[2:0]};
  ZLL_Main_compute410  instR48 (zll_main_compute410_inR4[5:3], zll_main_compute410_inR4[2:0], zll_main_compute410_outR4);
  assign zll_main_compute452_in = {zll_main_compute82_in[133:70], zll_main_compute82_in[69:6], zll_main_compute82_in[2:0], zll_main_compute82_in[5:3], zll_main_compute410_outR4};
  assign zll_main_compute173_in = {zll_main_compute452_in[136:73], zll_main_compute452_in[5:3], zll_main_compute452_in[2:0], 1'h0};
  assign zll_main_compute270_in = {zll_main_compute173_in[6:4], zll_main_compute173_in[3:1], 1'h0};
  ZLL_Main_compute270  instR49 (zll_main_compute270_in[6:4], zll_main_compute270_in[3:1], zll_main_compute270_in[0], zll_main_compute270_out);
  assign id_inR1 = {zll_main_compute173_in[3:1], zll_main_compute173_in[0]};
  assign zll_main_compute39_in = {zll_main_compute452_in[136:73], zll_main_compute452_in[72:9], zll_main_compute452_in[8:6], zll_main_compute452_in[5:3], (id_inR1[0] == 1'h1) ? id_inR1[3:1] : zll_main_compute270_out};
  assign zll_main_compute187_in = {zll_main_compute39_in[136:73], zll_main_compute39_in[2:0], zll_main_compute39_in[72:9], zll_main_compute39_in[8:6], zll_main_compute39_in[5:3], 3'h0};
  ZLL_Main_compute187  instR50 (zll_main_compute187_in[139:76], zll_main_compute187_in[75:73], zll_main_compute187_in[72:9], zll_main_compute187_in[8:6], zll_main_compute187_in[5:3], zll_main_compute187_in[2:0], zll_main_compute187_out);
  assign zll_main_compute187_inR1 = {zll_main_compute39_in[136:73], zll_main_compute39_in[2:0], zll_main_compute39_in[72:9], zll_main_compute39_in[8:6], zll_main_compute39_in[5:3], 3'h1};
  ZLL_Main_compute187  instR51 (zll_main_compute187_inR1[139:76], zll_main_compute187_inR1[75:73], zll_main_compute187_inR1[72:9], zll_main_compute187_inR1[8:6], zll_main_compute187_inR1[5:3], zll_main_compute187_inR1[2:0], zll_main_compute187_outR1);
  assign zll_main_compute187_inR2 = {zll_main_compute39_in[136:73], zll_main_compute39_in[2:0], zll_main_compute39_in[72:9], zll_main_compute39_in[8:6], zll_main_compute39_in[5:3], 3'h2};
  ZLL_Main_compute187  instR52 (zll_main_compute187_inR2[139:76], zll_main_compute187_inR2[75:73], zll_main_compute187_inR2[72:9], zll_main_compute187_inR2[8:6], zll_main_compute187_inR2[5:3], zll_main_compute187_inR2[2:0], zll_main_compute187_outR2);
  assign zll_main_compute187_inR3 = {zll_main_compute39_in[136:73], zll_main_compute39_in[2:0], zll_main_compute39_in[72:9], zll_main_compute39_in[8:6], zll_main_compute39_in[5:3], 3'h3};
  ZLL_Main_compute187  instR53 (zll_main_compute187_inR3[139:76], zll_main_compute187_inR3[75:73], zll_main_compute187_inR3[72:9], zll_main_compute187_inR3[8:6], zll_main_compute187_inR3[5:3], zll_main_compute187_inR3[2:0], zll_main_compute187_outR3);
  assign zll_main_compute187_inR4 = {zll_main_compute39_in[136:73], zll_main_compute39_in[2:0], zll_main_compute39_in[72:9], zll_main_compute39_in[8:6], zll_main_compute39_in[5:3], 3'h4};
  ZLL_Main_compute187  instR54 (zll_main_compute187_inR4[139:76], zll_main_compute187_inR4[75:73], zll_main_compute187_inR4[72:9], zll_main_compute187_inR4[8:6], zll_main_compute187_inR4[5:3], zll_main_compute187_inR4[2:0], zll_main_compute187_outR4);
  assign zll_main_compute187_inR5 = {zll_main_compute39_in[136:73], zll_main_compute39_in[2:0], zll_main_compute39_in[72:9], zll_main_compute39_in[8:6], zll_main_compute39_in[5:3], 3'h5};
  ZLL_Main_compute187  instR55 (zll_main_compute187_inR5[139:76], zll_main_compute187_inR5[75:73], zll_main_compute187_inR5[72:9], zll_main_compute187_inR5[8:6], zll_main_compute187_inR5[5:3], zll_main_compute187_inR5[2:0], zll_main_compute187_outR5);
  assign zll_main_compute187_inR6 = {zll_main_compute39_in[136:73], zll_main_compute39_in[2:0], zll_main_compute39_in[72:9], zll_main_compute39_in[8:6], zll_main_compute39_in[5:3], 3'h6};
  ZLL_Main_compute187  instR56 (zll_main_compute187_inR6[139:76], zll_main_compute187_inR6[75:73], zll_main_compute187_inR6[72:9], zll_main_compute187_inR6[8:6], zll_main_compute187_inR6[5:3], zll_main_compute187_inR6[2:0], zll_main_compute187_outR6);
  assign zll_main_compute187_inR7 = {zll_main_compute39_in[136:73], zll_main_compute39_in[2:0], zll_main_compute39_in[72:9], zll_main_compute39_in[8:6], zll_main_compute39_in[5:3], 3'h7};
  ZLL_Main_compute187  instR57 (zll_main_compute187_inR7[139:76], zll_main_compute187_inR7[75:73], zll_main_compute187_inR7[72:9], zll_main_compute187_inR7[8:6], zll_main_compute187_inR7[5:3], zll_main_compute187_inR7[2:0], zll_main_compute187_outR7);
  assign zll_main_compute258_in = {{zll_main_compute238_out, zll_main_compute238_outR1, zll_main_compute238_outR2, zll_main_compute238_outR3, zll_main_compute238_outR4, zll_main_compute238_outR5, zll_main_compute238_outR6, zll_main_compute238_outR7}, {zll_main_compute187_out, zll_main_compute187_outR1, zll_main_compute187_outR2, zll_main_compute187_outR3, zll_main_compute187_outR4, zll_main_compute187_outR5, zll_main_compute187_outR6, zll_main_compute187_outR7}};
  assign id_inR2 = zll_main_compute258_in[127:0];
  assign zll_main_loop2_in = {1'h0, {id_inR2[127:64], id_inR2[63:0]}};
  assign zll_main_loop_in = zll_main_loop2_in[128:0];
  assign {__padding, __out0, __out1} = {1'h1, zll_main_loop_in[127:0]};
endmodule

module ZLL_Main_compute439 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  output logic [0:0] res);
  logic [5:0] zll_main_compute235_in;
  logic [5:0] zll_main_compute377_in;
  logic [2:0] resize_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  assign zll_main_compute235_in = {arg0, arg1};
  assign zll_main_compute377_in = zll_main_compute235_in[5:0];
  assign resize_in = zll_main_compute377_in[5:3];
  assign resize_inR1 = zll_main_compute377_in[2:0];
  assign binop_in = {128'(resize_in[2:0]), 128'(resize_inR1[2:0])};
  assign res = binop_in[255:128] < binop_in[127:0];
endmodule

module ZLL_Main_compute412 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  input logic [63:0] arg2,
  output logic [7:0] res);
  logic [63:0] resize_in;
  logic [5:0] zll_main_compute368_in;
  logic [2:0] zll_main_compute368_out;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR2;
  assign resize_in = arg2;
  assign zll_main_compute368_in = {arg0, arg1};
  ZLL_Main_compute368  inst (zll_main_compute368_in[5:3], zll_main_compute368_in[2:0], zll_main_compute368_out);
  assign resize_inR1 = zll_main_compute368_out;
  assign binop_in = {128'h8, 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h8};
  assign binop_inR3 = {128'(resize_in[63:0]), binop_inR2[255:128] * binop_inR2[127:0]};
  assign resize_inR2 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign res = resize_inR2[7:0];
endmodule

module ZLL_Main_compute411 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  output logic [2:0] res);
  logic [5:0] zll_main_compute372_in;
  logic [5:0] zll_main_compute401_in;
  logic [2:0] resize_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR2;
  assign zll_main_compute372_in = {arg0, arg1};
  assign zll_main_compute401_in = zll_main_compute372_in[5:0];
  assign resize_in = zll_main_compute401_in[5:3];
  assign resize_inR1 = zll_main_compute401_in[2:0];
  assign binop_in = {128'(resize_in[2:0]), 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] + binop_in[127:0], 128'h8};
  assign resize_inR2 = binop_inR1[255:128] % binop_inR1[127:0];
  assign res = resize_inR2[2:0];
endmodule

module ZLL_Main_compute410 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  output logic [2:0] res);
  logic [5:0] zll_main_compute409_in;
  logic [5:0] zll_main_compute441_in;
  logic [2:0] resize_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR2;
  assign zll_main_compute409_in = {arg0, arg1};
  assign zll_main_compute441_in = zll_main_compute409_in[5:0];
  assign resize_in = zll_main_compute441_in[5:3];
  assign resize_inR1 = zll_main_compute441_in[2:0];
  assign binop_in = {128'(resize_in[2:0]), 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] / binop_in[127:0], 128'h8};
  assign resize_inR2 = binop_inR1[255:128] % binop_inR1[127:0];
  assign res = resize_inR2[2:0];
endmodule

module ZLL_Main_compute386 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  input logic [63:0] arg2,
  input logic [0:0] arg3,
  output logic [2:0] res);
  logic [6:0] zll_main_compute270_in;
  logic [2:0] zll_main_compute270_out;
  logic [3:0] id_in;
  assign zll_main_compute270_in = {arg0, arg1, 1'h0};
  ZLL_Main_compute270  inst (zll_main_compute270_in[6:4], zll_main_compute270_in[3:1], zll_main_compute270_in[0], zll_main_compute270_out);
  assign id_in = {arg1, arg3};
  assign res = (id_in[0] == 1'h1) ? id_in[3:1] : zll_main_compute270_out;
endmodule

module ZLL_Main_compute381 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  output logic [2:0] res);
  logic [5:0] zll_main_compute451_in;
  logic [5:0] zll_main_compute311_in;
  logic [2:0] resize_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR2;
  assign zll_main_compute451_in = {arg0, arg1};
  assign zll_main_compute311_in = zll_main_compute451_in[5:0];
  assign resize_in = zll_main_compute311_in[5:3];
  assign resize_inR1 = zll_main_compute311_in[2:0];
  assign binop_in = {128'(resize_in[2:0]), 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h8};
  assign resize_inR2 = binop_inR1[255:128] % binop_inR1[127:0];
  assign res = resize_inR2[2:0];
endmodule

module ZLL_Main_compute368 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  output logic [2:0] res);
  logic [5:0] zll_main_compute388_in;
  logic [5:0] zll_main_compute426_in;
  logic [2:0] resize_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR2;
  assign zll_main_compute388_in = {arg0, arg1};
  assign zll_main_compute426_in = zll_main_compute388_in[5:0];
  assign resize_in = zll_main_compute426_in[5:3];
  assign resize_inR1 = zll_main_compute426_in[2:0];
  assign binop_in = {128'(resize_in[2:0]), 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] * binop_in[127:0], 128'h8};
  assign resize_inR2 = binop_inR1[255:128] % binop_inR1[127:0];
  assign res = resize_inR2[2:0];
endmodule

module ZLL_Main_compute270 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  input logic [0:0] arg2,
  output logic [2:0] res);
  logic [6:0] zll_main_compute389_in;
  logic [5:0] zll_main_compute411_in;
  logic [2:0] zll_main_compute411_out;
  assign zll_main_compute389_in = {arg0, arg1, arg2};
  assign zll_main_compute411_in = {zll_main_compute389_in[3:1], zll_main_compute389_in[6:4]};
  ZLL_Main_compute411  inst (zll_main_compute411_in[5:3], zll_main_compute411_in[2:0], zll_main_compute411_out);
  assign res = zll_main_compute411_out;
endmodule

module ZLL_Main_compute238 (input logic [63:0] arg0,
  input logic [2:0] arg1,
  input logic [2:0] arg2,
  input logic [63:0] arg3,
  input logic [2:0] arg4,
  output logic [7:0] res);
  logic [2:0] zll_main_compute219_in;
  logic [0:0] zll_main_compute219_out;
  logic [137:0] zll_main_compute57_in;
  logic [2:0] zll_main_compute219_inR1;
  logic [0:0] zll_main_compute219_outR1;
  logic [73:0] zll_main_compute197_in;
  logic [73:0] zll_main_compute164_in;
  logic [63:0] resize_in;
  logic [5:0] zll_main_compute381_in;
  logic [2:0] zll_main_compute381_out;
  logic [5:0] zll_main_compute410_in;
  logic [2:0] zll_main_compute410_out;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR2;
  logic [70:0] zll_main_compute359_in;
  logic [63:0] resize_inR3;
  logic [5:0] zll_main_compute410_inR1;
  logic [2:0] zll_main_compute410_outR1;
  logic [2:0] resize_inR4;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR5;
  assign zll_main_compute219_in = arg4;
  ZLL_Main_compute219  inst (zll_main_compute219_in[2:0], zll_main_compute219_out);
  assign zll_main_compute57_in = {arg4, arg0, arg1, arg2, arg3, zll_main_compute219_out};
  assign zll_main_compute219_inR1 = zll_main_compute57_in[137:135];
  ZLL_Main_compute219  instR1 (zll_main_compute219_inR1[2:0], zll_main_compute219_outR1);
  assign zll_main_compute197_in = {zll_main_compute57_in[137:135], zll_main_compute57_in[70:68], zll_main_compute57_in[67:65], zll_main_compute57_in[64:1], zll_main_compute219_outR1};
  assign zll_main_compute164_in = {zll_main_compute197_in[73:71], zll_main_compute197_in[70:68], zll_main_compute197_in[67:65], zll_main_compute197_in[64:1], zll_main_compute197_in[0]};
  assign resize_in = zll_main_compute164_in[64:1];
  assign zll_main_compute381_in = {zll_main_compute164_in[73:71], zll_main_compute164_in[67:65]};
  ZLL_Main_compute381  instR2 (zll_main_compute381_in[5:3], zll_main_compute381_in[2:0], zll_main_compute381_out);
  assign zll_main_compute410_in = {zll_main_compute381_out, zll_main_compute164_in[70:68]};
  ZLL_Main_compute410  instR3 (zll_main_compute410_in[5:3], zll_main_compute410_in[2:0], zll_main_compute410_out);
  assign resize_inR1 = zll_main_compute410_out;
  assign binop_in = {128'h8, 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h8};
  assign binop_inR3 = {128'(resize_in[63:0]), binop_inR2[255:128] * binop_inR2[127:0]};
  assign resize_inR2 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign zll_main_compute359_in = {zll_main_compute57_in[137:135], zll_main_compute57_in[134:71], zll_main_compute57_in[70:68], zll_main_compute57_in[0]};
  assign resize_inR3 = zll_main_compute359_in[67:4];
  assign zll_main_compute410_inR1 = {zll_main_compute359_in[70:68], zll_main_compute359_in[3:1]};
  ZLL_Main_compute410  instR4 (zll_main_compute410_inR1[5:3], zll_main_compute410_inR1[2:0], zll_main_compute410_outR1);
  assign resize_inR4 = zll_main_compute410_outR1;
  assign binop_inR4 = {128'h8, 128'(resize_inR4[2:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h8};
  assign binop_inR7 = {128'(resize_inR3[63:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR5 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign res = (zll_main_compute359_in[0] == 1'h1) ? resize_inR5[7:0] : resize_inR2[7:0];
endmodule

module ZLL_Main_compute232 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  input logic [63:0] arg2,
  input logic [2:0] arg3,
  input logic [63:0] arg4,
  input logic [2:0] arg5,
  output logic [7:0] res);
  logic [5:0] zll_main_compute439_in;
  logic [0:0] zll_main_compute439_out;
  logic [140:0] zll_main_compute285_in;
  logic [5:0] zll_main_compute439_inR1;
  logic [0:0] zll_main_compute439_outR1;
  logic [76:0] zll_main_compute145_in;
  logic [76:0] zll_main_compute431_in;
  logic [63:0] resize_in;
  logic [5:0] zll_main_compute381_in;
  logic [2:0] zll_main_compute381_out;
  logic [5:0] zll_main_compute368_in;
  logic [2:0] zll_main_compute368_out;
  logic [5:0] zll_main_compute411_in;
  logic [2:0] zll_main_compute411_out;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR2;
  logic [73:0] zll_main_compute416_in;
  logic [63:0] resize_inR3;
  logic [5:0] zll_main_compute368_inR1;
  logic [2:0] zll_main_compute368_outR1;
  logic [5:0] zll_main_compute411_inR1;
  logic [2:0] zll_main_compute411_outR1;
  logic [2:0] resize_inR4;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR5;
  assign zll_main_compute439_in = {arg5, arg3};
  ZLL_Main_compute439  inst (zll_main_compute439_in[5:3], zll_main_compute439_in[2:0], zll_main_compute439_out);
  assign zll_main_compute285_in = {arg0, arg5, arg1, arg2, arg3, arg4, zll_main_compute439_out};
  assign zll_main_compute439_inR1 = {zll_main_compute285_in[137:135], zll_main_compute285_in[67:65]};
  ZLL_Main_compute439  instR1 (zll_main_compute439_inR1[5:3], zll_main_compute439_inR1[2:0], zll_main_compute439_outR1);
  assign zll_main_compute145_in = {zll_main_compute285_in[140:138], zll_main_compute285_in[137:135], zll_main_compute285_in[134:132], zll_main_compute285_in[67:65], zll_main_compute285_in[64:1], zll_main_compute439_outR1};
  assign zll_main_compute431_in = {zll_main_compute145_in[76:74], zll_main_compute145_in[73:71], zll_main_compute145_in[70:68], zll_main_compute145_in[67:65], zll_main_compute145_in[64:1], zll_main_compute145_in[0]};
  assign resize_in = zll_main_compute431_in[64:1];
  assign zll_main_compute381_in = {zll_main_compute431_in[73:71], zll_main_compute431_in[67:65]};
  ZLL_Main_compute381  instR2 (zll_main_compute381_in[5:3], zll_main_compute381_in[2:0], zll_main_compute381_out);
  assign zll_main_compute368_in = {zll_main_compute381_out, zll_main_compute431_in[70:68]};
  ZLL_Main_compute368  instR3 (zll_main_compute368_in[5:3], zll_main_compute368_in[2:0], zll_main_compute368_out);
  assign zll_main_compute411_in = {zll_main_compute368_out, zll_main_compute431_in[76:74]};
  ZLL_Main_compute411  instR4 (zll_main_compute411_in[5:3], zll_main_compute411_in[2:0], zll_main_compute411_out);
  assign resize_inR1 = zll_main_compute411_out;
  assign binop_in = {128'h8, 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h8};
  assign binop_inR3 = {128'(resize_in[63:0]), binop_inR2[255:128] * binop_inR2[127:0]};
  assign resize_inR2 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign zll_main_compute416_in = {zll_main_compute285_in[140:138], zll_main_compute285_in[137:135], zll_main_compute285_in[134:132], zll_main_compute285_in[131:68], zll_main_compute285_in[0]};
  assign resize_inR3 = zll_main_compute416_in[64:1];
  assign zll_main_compute368_inR1 = {zll_main_compute416_in[70:68], zll_main_compute416_in[67:65]};
  ZLL_Main_compute368  instR5 (zll_main_compute368_inR1[5:3], zll_main_compute368_inR1[2:0], zll_main_compute368_outR1);
  assign zll_main_compute411_inR1 = {zll_main_compute368_outR1, zll_main_compute416_in[73:71]};
  ZLL_Main_compute411  instR6 (zll_main_compute411_inR1[5:3], zll_main_compute411_inR1[2:0], zll_main_compute411_outR1);
  assign resize_inR4 = zll_main_compute411_outR1;
  assign binop_inR4 = {128'h8, 128'(resize_inR4[2:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h8};
  assign binop_inR7 = {128'(resize_inR3[63:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR5 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign res = (zll_main_compute416_in[0] == 1'h1) ? resize_inR5[7:0] : resize_inR2[7:0];
endmodule

module ZLL_Main_compute219 (input logic [2:0] arg0,
  output logic [0:0] res);
  logic [2:0] resize_in;
  logic [127:0] zll_main_compute366_in;
  logic [127:0] resize_inR1;
  logic [0:0] msbit_in;
  logic [0:0] rewire_prelude_not_in;
  logic [1:0] zll_rewire_prelude_not_in;
  logic [0:0] lit_in;
  assign resize_in = arg0;
  assign zll_main_compute366_in = 128'(resize_in[2:0]);
  assign resize_inR1 = zll_main_compute366_in[127:0];
  assign msbit_in = resize_inR1[0];
  assign rewire_prelude_not_in = msbit_in[0];
  assign zll_rewire_prelude_not_in = {rewire_prelude_not_in[0], rewire_prelude_not_in[0]};
  assign lit_in = zll_rewire_prelude_not_in[0];
  assign res = (lit_in[0] == 1'h1) ? 1'h0 : 1'h1;
endmodule

module ZLL_Main_compute215 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  input logic [63:0] arg2,
  input logic [63:0] arg3,
  input logic [2:0] arg4,
  input logic [2:0] arg5,
  output logic [7:0] res);
  logic [5:0] zll_main_compute439_in;
  logic [0:0] zll_main_compute439_out;
  logic [140:0] zll_main_compute81_in;
  logic [5:0] zll_main_compute439_inR1;
  logic [0:0] zll_main_compute439_outR1;
  logic [76:0] zll_main_compute37_in;
  logic [76:0] zll_main_compute162_in;
  logic [63:0] resize_in;
  logic [5:0] zll_main_compute381_in;
  logic [2:0] zll_main_compute381_out;
  logic [5:0] zll_main_compute368_in;
  logic [2:0] zll_main_compute368_out;
  logic [5:0] zll_main_compute411_in;
  logic [2:0] zll_main_compute411_out;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR2;
  logic [73:0] zll_main_compute230_in;
  logic [63:0] resize_inR3;
  logic [5:0] zll_main_compute368_inR1;
  logic [2:0] zll_main_compute368_outR1;
  logic [5:0] zll_main_compute411_inR1;
  logic [2:0] zll_main_compute411_outR1;
  logic [2:0] resize_inR4;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR5;
  assign zll_main_compute439_in = {arg5, arg4};
  ZLL_Main_compute439  inst (zll_main_compute439_in[5:3], zll_main_compute439_in[2:0], zll_main_compute439_out);
  assign zll_main_compute81_in = {arg0, arg1, arg2, arg3, arg4, arg5, zll_main_compute439_out};
  assign zll_main_compute439_inR1 = {zll_main_compute81_in[3:1], zll_main_compute81_in[6:4]};
  ZLL_Main_compute439  instR1 (zll_main_compute439_inR1[5:3], zll_main_compute439_inR1[2:0], zll_main_compute439_outR1);
  assign zll_main_compute37_in = {zll_main_compute81_in[140:138], zll_main_compute81_in[137:135], zll_main_compute81_in[70:7], zll_main_compute81_in[6:4], zll_main_compute81_in[3:1], zll_main_compute439_outR1};
  assign zll_main_compute162_in = {zll_main_compute37_in[76:74], zll_main_compute37_in[73:71], zll_main_compute37_in[70:7], zll_main_compute37_in[6:4], zll_main_compute37_in[3:1], zll_main_compute37_in[0]};
  assign resize_in = zll_main_compute162_in[70:7];
  assign zll_main_compute381_in = {zll_main_compute162_in[3:1], zll_main_compute162_in[6:4]};
  ZLL_Main_compute381  instR2 (zll_main_compute381_in[5:3], zll_main_compute381_in[2:0], zll_main_compute381_out);
  assign zll_main_compute368_in = {zll_main_compute381_out, zll_main_compute162_in[76:74]};
  ZLL_Main_compute368  instR3 (zll_main_compute368_in[5:3], zll_main_compute368_in[2:0], zll_main_compute368_out);
  assign zll_main_compute411_in = {zll_main_compute368_out, zll_main_compute162_in[73:71]};
  ZLL_Main_compute411  instR4 (zll_main_compute411_in[5:3], zll_main_compute411_in[2:0], zll_main_compute411_out);
  assign resize_inR1 = zll_main_compute411_out;
  assign binop_in = {128'h8, 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h8};
  assign binop_inR3 = {128'(resize_in[63:0]), binop_inR2[255:128] * binop_inR2[127:0]};
  assign resize_inR2 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign zll_main_compute230_in = {zll_main_compute81_in[140:138], zll_main_compute81_in[137:135], zll_main_compute81_in[134:71], zll_main_compute81_in[3:1], zll_main_compute81_in[0]};
  assign resize_inR3 = zll_main_compute230_in[67:4];
  assign zll_main_compute368_inR1 = {zll_main_compute230_in[3:1], zll_main_compute230_in[73:71]};
  ZLL_Main_compute368  instR5 (zll_main_compute368_inR1[5:3], zll_main_compute368_inR1[2:0], zll_main_compute368_outR1);
  assign zll_main_compute411_inR1 = {zll_main_compute368_outR1, zll_main_compute230_in[70:68]};
  ZLL_Main_compute411  instR6 (zll_main_compute411_inR1[5:3], zll_main_compute411_inR1[2:0], zll_main_compute411_outR1);
  assign resize_inR4 = zll_main_compute411_outR1;
  assign binop_inR4 = {128'h8, 128'(resize_inR4[2:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h8};
  assign binop_inR7 = {128'(resize_inR3[63:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR5 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign res = (zll_main_compute230_in[0] == 1'h1) ? resize_inR5[7:0] : resize_inR2[7:0];
endmodule

module ZLL_Main_compute187 (input logic [63:0] arg0,
  input logic [2:0] arg1,
  input logic [63:0] arg2,
  input logic [2:0] arg3,
  input logic [2:0] arg4,
  input logic [2:0] arg5,
  output logic [7:0] res);
  logic [2:0] zll_main_compute219_in;
  logic [0:0] zll_main_compute219_out;
  logic [140:0] zll_main_compute131_in;
  logic [2:0] zll_main_compute219_inR1;
  logic [0:0] zll_main_compute219_outR1;
  logic [76:0] zll_main_compute298_in;
  logic [76:0] zll_main_compute338_in;
  logic [63:0] resize_in;
  logic [5:0] zll_main_compute381_in;
  logic [2:0] zll_main_compute381_out;
  logic [5:0] zll_main_compute410_in;
  logic [2:0] zll_main_compute410_out;
  logic [5:0] zll_main_compute411_in;
  logic [2:0] zll_main_compute411_out;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR2;
  logic [73:0] zll_main_compute76_in;
  logic [63:0] resize_inR3;
  logic [5:0] zll_main_compute410_inR1;
  logic [2:0] zll_main_compute410_outR1;
  logic [5:0] zll_main_compute411_inR1;
  logic [2:0] zll_main_compute411_outR1;
  logic [2:0] resize_inR4;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR5;
  assign zll_main_compute219_in = arg5;
  ZLL_Main_compute219  inst (zll_main_compute219_in[2:0], zll_main_compute219_out);
  assign zll_main_compute131_in = {arg0, arg1, arg2, arg3, arg5, arg4, zll_main_compute219_out};
  assign zll_main_compute219_inR1 = zll_main_compute131_in[6:4];
  ZLL_Main_compute219  instR1 (zll_main_compute219_inR1[2:0], zll_main_compute219_outR1);
  assign zll_main_compute298_in = {zll_main_compute131_in[76:74], zll_main_compute131_in[73:10], zll_main_compute131_in[9:7], zll_main_compute131_in[6:4], zll_main_compute131_in[3:1], zll_main_compute219_outR1};
  assign zll_main_compute338_in = {zll_main_compute298_in[76:74], zll_main_compute298_in[73:10], zll_main_compute298_in[9:7], zll_main_compute298_in[6:4], zll_main_compute298_in[3:1], zll_main_compute298_in[0]};
  assign resize_in = zll_main_compute338_in[73:10];
  assign zll_main_compute381_in = {zll_main_compute338_in[6:4], zll_main_compute338_in[3:1]};
  ZLL_Main_compute381  instR2 (zll_main_compute381_in[5:3], zll_main_compute381_in[2:0], zll_main_compute381_out);
  assign zll_main_compute410_in = {zll_main_compute381_out, zll_main_compute338_in[9:7]};
  ZLL_Main_compute410  instR3 (zll_main_compute410_in[5:3], zll_main_compute410_in[2:0], zll_main_compute410_out);
  assign zll_main_compute411_in = {zll_main_compute338_in[76:74], zll_main_compute410_out};
  ZLL_Main_compute411  instR4 (zll_main_compute411_in[5:3], zll_main_compute411_in[2:0], zll_main_compute411_out);
  assign resize_inR1 = zll_main_compute411_out;
  assign binop_in = {128'h8, 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h8};
  assign binop_inR3 = {128'(resize_in[63:0]), binop_inR2[255:128] * binop_inR2[127:0]};
  assign resize_inR2 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign zll_main_compute76_in = {zll_main_compute131_in[140:77], zll_main_compute131_in[76:74], zll_main_compute131_in[9:7], zll_main_compute131_in[6:4], zll_main_compute131_in[0]};
  assign resize_inR3 = zll_main_compute76_in[73:10];
  assign zll_main_compute410_inR1 = {zll_main_compute76_in[3:1], zll_main_compute76_in[6:4]};
  ZLL_Main_compute410  instR5 (zll_main_compute410_inR1[5:3], zll_main_compute410_inR1[2:0], zll_main_compute410_outR1);
  assign zll_main_compute411_inR1 = {zll_main_compute76_in[9:7], zll_main_compute410_outR1};
  ZLL_Main_compute411  instR6 (zll_main_compute411_inR1[5:3], zll_main_compute411_inR1[2:0], zll_main_compute411_outR1);
  assign resize_inR4 = zll_main_compute411_outR1;
  assign binop_inR4 = {128'h8, 128'(resize_inR4[2:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h8};
  assign binop_inR7 = {128'(resize_inR3[63:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR5 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign res = (zll_main_compute76_in[0] == 1'h1) ? resize_inR5[7:0] : resize_inR2[7:0];
endmodule

module ZLL_Main_compute126 (input logic [2:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  input logic [63:0] arg3,
  input logic [2:0] arg4,
  output logic [7:0] res);
  logic [5:0] zll_main_compute439_in;
  logic [0:0] zll_main_compute439_out;
  logic [137:0] zll_main_compute139_in;
  logic [5:0] zll_main_compute439_inR1;
  logic [0:0] zll_main_compute439_outR1;
  logic [73:0] zll_main_compute402_in;
  logic [73:0] zll_main_compute133_in;
  logic [63:0] resize_in;
  logic [5:0] zll_main_compute381_in;
  logic [2:0] zll_main_compute381_out;
  logic [5:0] zll_main_compute368_in;
  logic [2:0] zll_main_compute368_out;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR2;
  logic [70:0] zll_main_compute412_in;
  logic [7:0] zll_main_compute412_out;
  assign zll_main_compute439_in = {arg4, arg2};
  ZLL_Main_compute439  inst (zll_main_compute439_in[5:3], zll_main_compute439_in[2:0], zll_main_compute439_out);
  assign zll_main_compute139_in = {arg4, arg0, arg1, arg2, arg3, zll_main_compute439_out};
  assign zll_main_compute439_inR1 = {zll_main_compute139_in[137:135], zll_main_compute139_in[67:65]};
  ZLL_Main_compute439  instR1 (zll_main_compute439_inR1[5:3], zll_main_compute439_inR1[2:0], zll_main_compute439_outR1);
  assign zll_main_compute402_in = {zll_main_compute139_in[137:135], zll_main_compute139_in[134:132], zll_main_compute139_in[67:65], zll_main_compute139_in[64:1], zll_main_compute439_outR1};
  assign zll_main_compute133_in = {zll_main_compute402_in[73:71], zll_main_compute402_in[70:68], zll_main_compute402_in[67:65], zll_main_compute402_in[64:1], zll_main_compute402_in[0]};
  assign resize_in = zll_main_compute133_in[64:1];
  assign zll_main_compute381_in = {zll_main_compute133_in[73:71], zll_main_compute133_in[67:65]};
  ZLL_Main_compute381  instR2 (zll_main_compute381_in[5:3], zll_main_compute381_in[2:0], zll_main_compute381_out);
  assign zll_main_compute368_in = {zll_main_compute381_out, zll_main_compute133_in[70:68]};
  ZLL_Main_compute368  instR3 (zll_main_compute368_in[5:3], zll_main_compute368_in[2:0], zll_main_compute368_out);
  assign resize_inR1 = zll_main_compute368_out;
  assign binop_in = {128'h8, 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h8};
  assign binop_inR3 = {128'(resize_in[63:0]), binop_inR2[255:128] * binop_inR2[127:0]};
  assign resize_inR2 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign zll_main_compute412_in = {zll_main_compute139_in[137:135], zll_main_compute139_in[134:132], zll_main_compute139_in[131:68], zll_main_compute139_in[0]};
  ZLL_Main_compute412  instR4 (zll_main_compute412_in[70:68], zll_main_compute412_in[67:65], zll_main_compute412_in[64:1], zll_main_compute412_out);
  assign res = (zll_main_compute412_in[0] == 1'h1) ? zll_main_compute412_out : resize_inR2[7:0];
endmodule

module ZLL_Main_compute41 (input logic [2:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  input logic [63:0] arg3,
  input logic [2:0] arg4,
  output logic [7:0] res);
  logic [5:0] zll_main_compute439_in;
  logic [0:0] zll_main_compute439_out;
  logic [137:0] zll_main_compute357_in;
  logic [5:0] zll_main_compute439_inR1;
  logic [0:0] zll_main_compute439_outR1;
  logic [73:0] zll_main_compute80_in;
  logic [73:0] zll_main_compute251_in;
  logic [63:0] resize_in;
  logic [5:0] zll_main_compute381_in;
  logic [2:0] zll_main_compute381_out;
  logic [5:0] zll_main_compute368_in;
  logic [2:0] zll_main_compute368_out;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR2;
  logic [70:0] zll_main_compute412_in;
  logic [7:0] zll_main_compute412_out;
  assign zll_main_compute439_in = {arg4, arg2};
  ZLL_Main_compute439  inst (zll_main_compute439_in[5:3], zll_main_compute439_in[2:0], zll_main_compute439_out);
  assign zll_main_compute357_in = {arg4, arg0, arg1, arg2, arg3, zll_main_compute439_out};
  assign zll_main_compute439_inR1 = {zll_main_compute357_in[137:135], zll_main_compute357_in[67:65]};
  ZLL_Main_compute439  instR1 (zll_main_compute439_inR1[5:3], zll_main_compute439_inR1[2:0], zll_main_compute439_outR1);
  assign zll_main_compute80_in = {zll_main_compute357_in[137:135], zll_main_compute357_in[134:132], zll_main_compute357_in[131:68], zll_main_compute357_in[67:65], zll_main_compute439_outR1};
  assign zll_main_compute251_in = {zll_main_compute80_in[73:71], zll_main_compute80_in[70:68], zll_main_compute80_in[67:4], zll_main_compute80_in[3:1], zll_main_compute80_in[0]};
  assign resize_in = zll_main_compute251_in[67:4];
  assign zll_main_compute381_in = {zll_main_compute251_in[73:71], zll_main_compute251_in[3:1]};
  ZLL_Main_compute381  instR2 (zll_main_compute381_in[5:3], zll_main_compute381_in[2:0], zll_main_compute381_out);
  assign zll_main_compute368_in = {zll_main_compute381_out, zll_main_compute251_in[70:68]};
  ZLL_Main_compute368  instR3 (zll_main_compute368_in[5:3], zll_main_compute368_in[2:0], zll_main_compute368_out);
  assign resize_inR1 = zll_main_compute368_out;
  assign binop_in = {128'h8, 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h8};
  assign binop_inR3 = {128'(resize_in[63:0]), binop_inR2[255:128] * binop_inR2[127:0]};
  assign resize_inR2 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign zll_main_compute412_in = {zll_main_compute357_in[137:135], zll_main_compute357_in[134:132], zll_main_compute357_in[64:1], zll_main_compute357_in[0]};
  ZLL_Main_compute412  instR4 (zll_main_compute412_in[70:68], zll_main_compute412_in[67:65], zll_main_compute412_in[64:1], zll_main_compute412_out);
  assign res = (zll_main_compute412_in[0] == 1'h1) ? zll_main_compute412_out : resize_inR2[7:0];
endmodule