module top_level (input logic [1:0] __in0,
  output logic [1:0] __out0);
  logic [0:0] __continue;
  assign {__continue, __out0} = 2'h1;
endmodule