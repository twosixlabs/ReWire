module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [99:0] __in0,
  output logic [99:0] __out0,
  output logic [99:0] __out1,
  output logic [99:0] __out2,
  output logic [99:0] __out3);
  logic [100:0] gzdLLzicase11834;
  logic [401:0] callRes;
  logic [100:0] gzdLLzicase11834R1;
  logic [401:0] callResR1;
  logic [0:0] __continue;
  logic [0:0] __resumption_tag;
  logic [0:0] __resumption_tag_next;
  assign gzdLLzicase11834 = {__resumption_tag, __in0};
  zdLLzicase11834  zdLLzicase11834 (gzdLLzicase11834[99:0], callRes);
  assign gzdLLzicase11834R1 = {__resumption_tag, __in0};
  zdLLzicase11834  zdLLzicase11834R1 (gzdLLzicase11834R1[99:0], callResR1);
  assign {__continue, __out0, __out1, __out2, __out3, __resumption_tag_next} = (gzdLLzicase11834R1[100] == 1'h0) ? callResR1 : callRes;
  initial __resumption_tag <= 1'h1;
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      __resumption_tag <= 1'h1;
    end else begin
      __resumption_tag <= __resumption_tag_next;
    end
  end
endmodule

module zdLLzicase11834 (input logic [99:0] arg0,
  output logic [401:0] res);
  logic [99:0] gMainzidev;
  logic [106:0] gzdLLzilambda11768;
  logic [0:0] callRes;
  logic [106:0] gzdLLzilambda11768R1;
  logic [0:0] callResR1;
  logic [106:0] gzdLLzilambda11768R2;
  logic [0:0] callResR2;
  logic [106:0] gzdLLzilambda11768R3;
  logic [0:0] callResR3;
  logic [106:0] gzdLLzilambda11768R4;
  logic [0:0] callResR4;
  logic [106:0] gzdLLzilambda11768R5;
  logic [0:0] callResR5;
  logic [106:0] gzdLLzilambda11768R6;
  logic [0:0] callResR6;
  logic [106:0] gzdLLzilambda11768R7;
  logic [0:0] callResR7;
  logic [106:0] gzdLLzilambda11768R8;
  logic [0:0] callResR8;
  logic [106:0] gzdLLzilambda11768R9;
  logic [0:0] callResR9;
  logic [106:0] gzdLLzilambda11768R10;
  logic [0:0] callResR10;
  logic [106:0] gzdLLzilambda11768R11;
  logic [0:0] callResR11;
  logic [106:0] gzdLLzilambda11768R12;
  logic [0:0] callResR12;
  logic [106:0] gzdLLzilambda11768R13;
  logic [0:0] callResR13;
  logic [106:0] gzdLLzilambda11768R14;
  logic [0:0] callResR14;
  logic [106:0] gzdLLzilambda11768R15;
  logic [0:0] callResR15;
  logic [106:0] gzdLLzilambda11768R16;
  logic [0:0] callResR16;
  logic [106:0] gzdLLzilambda11768R17;
  logic [0:0] callResR17;
  logic [106:0] gzdLLzilambda11768R18;
  logic [0:0] callResR18;
  logic [106:0] gzdLLzilambda11768R19;
  logic [0:0] callResR19;
  logic [106:0] gzdLLzilambda11768R20;
  logic [0:0] callResR20;
  logic [106:0] gzdLLzilambda11768R21;
  logic [0:0] callResR21;
  logic [106:0] gzdLLzilambda11768R22;
  logic [0:0] callResR22;
  logic [106:0] gzdLLzilambda11768R23;
  logic [0:0] callResR23;
  logic [106:0] gzdLLzilambda11768R24;
  logic [0:0] callResR24;
  logic [106:0] gzdLLzilambda11768R25;
  logic [0:0] callResR25;
  logic [106:0] gzdLLzilambda11768R26;
  logic [0:0] callResR26;
  logic [106:0] gzdLLzilambda11768R27;
  logic [0:0] callResR27;
  logic [106:0] gzdLLzilambda11768R28;
  logic [0:0] callResR28;
  logic [106:0] gzdLLzilambda11768R29;
  logic [0:0] callResR29;
  logic [106:0] gzdLLzilambda11768R30;
  logic [0:0] callResR30;
  logic [106:0] gzdLLzilambda11768R31;
  logic [0:0] callResR31;
  logic [106:0] gzdLLzilambda11768R32;
  logic [0:0] callResR32;
  logic [106:0] gzdLLzilambda11768R33;
  logic [0:0] callResR33;
  logic [106:0] gzdLLzilambda11768R34;
  logic [0:0] callResR34;
  logic [106:0] gzdLLzilambda11768R35;
  logic [0:0] callResR35;
  logic [106:0] gzdLLzilambda11768R36;
  logic [0:0] callResR36;
  logic [106:0] gzdLLzilambda11768R37;
  logic [0:0] callResR37;
  logic [106:0] gzdLLzilambda11768R38;
  logic [0:0] callResR38;
  logic [106:0] gzdLLzilambda11768R39;
  logic [0:0] callResR39;
  logic [106:0] gzdLLzilambda11768R40;
  logic [0:0] callResR40;
  logic [106:0] gzdLLzilambda11768R41;
  logic [0:0] callResR41;
  logic [106:0] gzdLLzilambda11768R42;
  logic [0:0] callResR42;
  logic [106:0] gzdLLzilambda11768R43;
  logic [0:0] callResR43;
  logic [106:0] gzdLLzilambda11768R44;
  logic [0:0] callResR44;
  logic [106:0] gzdLLzilambda11768R45;
  logic [0:0] callResR45;
  logic [106:0] gzdLLzilambda11768R46;
  logic [0:0] callResR46;
  logic [106:0] gzdLLzilambda11768R47;
  logic [0:0] callResR47;
  logic [106:0] gzdLLzilambda11768R48;
  logic [0:0] callResR48;
  logic [106:0] gzdLLzilambda11768R49;
  logic [0:0] callResR49;
  logic [106:0] gzdLLzilambda11768R50;
  logic [0:0] callResR50;
  logic [106:0] gzdLLzilambda11768R51;
  logic [0:0] callResR51;
  logic [106:0] gzdLLzilambda11768R52;
  logic [0:0] callResR52;
  logic [106:0] gzdLLzilambda11768R53;
  logic [0:0] callResR53;
  logic [106:0] gzdLLzilambda11768R54;
  logic [0:0] callResR54;
  logic [106:0] gzdLLzilambda11768R55;
  logic [0:0] callResR55;
  logic [106:0] gzdLLzilambda11768R56;
  logic [0:0] callResR56;
  logic [106:0] gzdLLzilambda11768R57;
  logic [0:0] callResR57;
  logic [106:0] gzdLLzilambda11768R58;
  logic [0:0] callResR58;
  logic [106:0] gzdLLzilambda11768R59;
  logic [0:0] callResR59;
  logic [106:0] gzdLLzilambda11768R60;
  logic [0:0] callResR60;
  logic [106:0] gzdLLzilambda11768R61;
  logic [0:0] callResR61;
  logic [106:0] gzdLLzilambda11768R62;
  logic [0:0] callResR62;
  logic [106:0] gzdLLzilambda11768R63;
  logic [0:0] callResR63;
  logic [106:0] gzdLLzilambda11768R64;
  logic [0:0] callResR64;
  logic [106:0] gzdLLzilambda11768R65;
  logic [0:0] callResR65;
  logic [106:0] gzdLLzilambda11768R66;
  logic [0:0] callResR66;
  logic [106:0] gzdLLzilambda11768R67;
  logic [0:0] callResR67;
  logic [106:0] gzdLLzilambda11768R68;
  logic [0:0] callResR68;
  logic [106:0] gzdLLzilambda11768R69;
  logic [0:0] callResR69;
  logic [106:0] gzdLLzilambda11768R70;
  logic [0:0] callResR70;
  logic [106:0] gzdLLzilambda11768R71;
  logic [0:0] callResR71;
  logic [106:0] gzdLLzilambda11768R72;
  logic [0:0] callResR72;
  logic [106:0] gzdLLzilambda11768R73;
  logic [0:0] callResR73;
  logic [106:0] gzdLLzilambda11768R74;
  logic [0:0] callResR74;
  logic [106:0] gzdLLzilambda11768R75;
  logic [0:0] callResR75;
  logic [106:0] gzdLLzilambda11768R76;
  logic [0:0] callResR76;
  logic [106:0] gzdLLzilambda11768R77;
  logic [0:0] callResR77;
  logic [106:0] gzdLLzilambda11768R78;
  logic [0:0] callResR78;
  logic [106:0] gzdLLzilambda11768R79;
  logic [0:0] callResR79;
  logic [106:0] gzdLLzilambda11768R80;
  logic [0:0] callResR80;
  logic [106:0] gzdLLzilambda11768R81;
  logic [0:0] callResR81;
  logic [106:0] gzdLLzilambda11768R82;
  logic [0:0] callResR82;
  logic [106:0] gzdLLzilambda11768R83;
  logic [0:0] callResR83;
  logic [106:0] gzdLLzilambda11768R84;
  logic [0:0] callResR84;
  logic [106:0] gzdLLzilambda11768R85;
  logic [0:0] callResR85;
  logic [106:0] gzdLLzilambda11768R86;
  logic [0:0] callResR86;
  logic [106:0] gzdLLzilambda11768R87;
  logic [0:0] callResR87;
  logic [106:0] gzdLLzilambda11768R88;
  logic [0:0] callResR88;
  logic [106:0] gzdLLzilambda11768R89;
  logic [0:0] callResR89;
  logic [106:0] gzdLLzilambda11768R90;
  logic [0:0] callResR90;
  logic [106:0] gzdLLzilambda11768R91;
  logic [0:0] callResR91;
  logic [106:0] gzdLLzilambda11768R92;
  logic [0:0] callResR92;
  logic [106:0] gzdLLzilambda11768R93;
  logic [0:0] callResR93;
  logic [106:0] gzdLLzilambda11768R94;
  logic [0:0] callResR94;
  logic [106:0] gzdLLzilambda11768R95;
  logic [0:0] callResR95;
  logic [106:0] gzdLLzilambda11768R96;
  logic [0:0] callResR96;
  logic [106:0] gzdLLzilambda11768R97;
  logic [0:0] callResR97;
  logic [106:0] gzdLLzilambda11768R98;
  logic [0:0] callResR98;
  logic [106:0] gzdLLzilambda11768R99;
  logic [0:0] callResR99;
  logic [106:0] gzdLLzilambda11777;
  logic [0:0] callResR100;
  logic [106:0] gzdLLzilambda11777R1;
  logic [0:0] callResR101;
  logic [106:0] gzdLLzilambda11777R2;
  logic [0:0] callResR102;
  logic [106:0] gzdLLzilambda11777R3;
  logic [0:0] callResR103;
  logic [106:0] gzdLLzilambda11777R4;
  logic [0:0] callResR104;
  logic [106:0] gzdLLzilambda11777R5;
  logic [0:0] callResR105;
  logic [106:0] gzdLLzilambda11777R6;
  logic [0:0] callResR106;
  logic [106:0] gzdLLzilambda11777R7;
  logic [0:0] callResR107;
  logic [106:0] gzdLLzilambda11777R8;
  logic [0:0] callResR108;
  logic [106:0] gzdLLzilambda11777R9;
  logic [0:0] callResR109;
  logic [106:0] gzdLLzilambda11777R10;
  logic [0:0] callResR110;
  logic [106:0] gzdLLzilambda11777R11;
  logic [0:0] callResR111;
  logic [106:0] gzdLLzilambda11777R12;
  logic [0:0] callResR112;
  logic [106:0] gzdLLzilambda11777R13;
  logic [0:0] callResR113;
  logic [106:0] gzdLLzilambda11777R14;
  logic [0:0] callResR114;
  logic [106:0] gzdLLzilambda11777R15;
  logic [0:0] callResR115;
  logic [106:0] gzdLLzilambda11777R16;
  logic [0:0] callResR116;
  logic [106:0] gzdLLzilambda11777R17;
  logic [0:0] callResR117;
  logic [106:0] gzdLLzilambda11777R18;
  logic [0:0] callResR118;
  logic [106:0] gzdLLzilambda11777R19;
  logic [0:0] callResR119;
  logic [106:0] gzdLLzilambda11777R20;
  logic [0:0] callResR120;
  logic [106:0] gzdLLzilambda11777R21;
  logic [0:0] callResR121;
  logic [106:0] gzdLLzilambda11777R22;
  logic [0:0] callResR122;
  logic [106:0] gzdLLzilambda11777R23;
  logic [0:0] callResR123;
  logic [106:0] gzdLLzilambda11777R24;
  logic [0:0] callResR124;
  logic [106:0] gzdLLzilambda11777R25;
  logic [0:0] callResR125;
  logic [106:0] gzdLLzilambda11777R26;
  logic [0:0] callResR126;
  logic [106:0] gzdLLzilambda11777R27;
  logic [0:0] callResR127;
  logic [106:0] gzdLLzilambda11777R28;
  logic [0:0] callResR128;
  logic [106:0] gzdLLzilambda11777R29;
  logic [0:0] callResR129;
  logic [106:0] gzdLLzilambda11777R30;
  logic [0:0] callResR130;
  logic [106:0] gzdLLzilambda11777R31;
  logic [0:0] callResR131;
  logic [106:0] gzdLLzilambda11777R32;
  logic [0:0] callResR132;
  logic [106:0] gzdLLzilambda11777R33;
  logic [0:0] callResR133;
  logic [106:0] gzdLLzilambda11777R34;
  logic [0:0] callResR134;
  logic [106:0] gzdLLzilambda11777R35;
  logic [0:0] callResR135;
  logic [106:0] gzdLLzilambda11777R36;
  logic [0:0] callResR136;
  logic [106:0] gzdLLzilambda11777R37;
  logic [0:0] callResR137;
  logic [106:0] gzdLLzilambda11777R38;
  logic [0:0] callResR138;
  logic [106:0] gzdLLzilambda11777R39;
  logic [0:0] callResR139;
  logic [106:0] gzdLLzilambda11777R40;
  logic [0:0] callResR140;
  logic [106:0] gzdLLzilambda11777R41;
  logic [0:0] callResR141;
  logic [106:0] gzdLLzilambda11777R42;
  logic [0:0] callResR142;
  logic [106:0] gzdLLzilambda11777R43;
  logic [0:0] callResR143;
  logic [106:0] gzdLLzilambda11777R44;
  logic [0:0] callResR144;
  logic [106:0] gzdLLzilambda11777R45;
  logic [0:0] callResR145;
  logic [106:0] gzdLLzilambda11777R46;
  logic [0:0] callResR146;
  logic [106:0] gzdLLzilambda11777R47;
  logic [0:0] callResR147;
  logic [106:0] gzdLLzilambda11777R48;
  logic [0:0] callResR148;
  logic [106:0] gzdLLzilambda11777R49;
  logic [0:0] callResR149;
  logic [106:0] gzdLLzilambda11777R50;
  logic [0:0] callResR150;
  logic [106:0] gzdLLzilambda11777R51;
  logic [0:0] callResR151;
  logic [106:0] gzdLLzilambda11777R52;
  logic [0:0] callResR152;
  logic [106:0] gzdLLzilambda11777R53;
  logic [0:0] callResR153;
  logic [106:0] gzdLLzilambda11777R54;
  logic [0:0] callResR154;
  logic [106:0] gzdLLzilambda11777R55;
  logic [0:0] callResR155;
  logic [106:0] gzdLLzilambda11777R56;
  logic [0:0] callResR156;
  logic [106:0] gzdLLzilambda11777R57;
  logic [0:0] callResR157;
  logic [106:0] gzdLLzilambda11777R58;
  logic [0:0] callResR158;
  logic [106:0] gzdLLzilambda11777R59;
  logic [0:0] callResR159;
  logic [106:0] gzdLLzilambda11777R60;
  logic [0:0] callResR160;
  logic [106:0] gzdLLzilambda11777R61;
  logic [0:0] callResR161;
  logic [106:0] gzdLLzilambda11777R62;
  logic [0:0] callResR162;
  logic [106:0] gzdLLzilambda11777R63;
  logic [0:0] callResR163;
  logic [106:0] gzdLLzilambda11777R64;
  logic [0:0] callResR164;
  logic [106:0] gzdLLzilambda11777R65;
  logic [0:0] callResR165;
  logic [106:0] gzdLLzilambda11777R66;
  logic [0:0] callResR166;
  logic [106:0] gzdLLzilambda11777R67;
  logic [0:0] callResR167;
  logic [106:0] gzdLLzilambda11777R68;
  logic [0:0] callResR168;
  logic [106:0] gzdLLzilambda11777R69;
  logic [0:0] callResR169;
  logic [106:0] gzdLLzilambda11777R70;
  logic [0:0] callResR170;
  logic [106:0] gzdLLzilambda11777R71;
  logic [0:0] callResR171;
  logic [106:0] gzdLLzilambda11777R72;
  logic [0:0] callResR172;
  logic [106:0] gzdLLzilambda11777R73;
  logic [0:0] callResR173;
  logic [106:0] gzdLLzilambda11777R74;
  logic [0:0] callResR174;
  logic [106:0] gzdLLzilambda11777R75;
  logic [0:0] callResR175;
  logic [106:0] gzdLLzilambda11777R76;
  logic [0:0] callResR176;
  logic [106:0] gzdLLzilambda11777R77;
  logic [0:0] callResR177;
  logic [106:0] gzdLLzilambda11777R78;
  logic [0:0] callResR178;
  logic [106:0] gzdLLzilambda11777R79;
  logic [0:0] callResR179;
  logic [106:0] gzdLLzilambda11777R80;
  logic [0:0] callResR180;
  logic [106:0] gzdLLzilambda11777R81;
  logic [0:0] callResR181;
  logic [106:0] gzdLLzilambda11777R82;
  logic [0:0] callResR182;
  logic [106:0] gzdLLzilambda11777R83;
  logic [0:0] callResR183;
  logic [106:0] gzdLLzilambda11777R84;
  logic [0:0] callResR184;
  logic [106:0] gzdLLzilambda11777R85;
  logic [0:0] callResR185;
  logic [106:0] gzdLLzilambda11777R86;
  logic [0:0] callResR186;
  logic [106:0] gzdLLzilambda11777R87;
  logic [0:0] callResR187;
  logic [106:0] gzdLLzilambda11777R88;
  logic [0:0] callResR188;
  logic [106:0] gzdLLzilambda11777R89;
  logic [0:0] callResR189;
  logic [106:0] gzdLLzilambda11777R90;
  logic [0:0] callResR190;
  logic [106:0] gzdLLzilambda11777R91;
  logic [0:0] callResR191;
  logic [106:0] gzdLLzilambda11777R92;
  logic [0:0] callResR192;
  logic [106:0] gzdLLzilambda11777R93;
  logic [0:0] callResR193;
  logic [106:0] gzdLLzilambda11777R94;
  logic [0:0] callResR194;
  logic [106:0] gzdLLzilambda11777R95;
  logic [0:0] callResR195;
  logic [106:0] gzdLLzilambda11777R96;
  logic [0:0] callResR196;
  logic [106:0] gzdLLzilambda11777R97;
  logic [0:0] callResR197;
  logic [106:0] gzdLLzilambda11777R98;
  logic [0:0] callResR198;
  logic [106:0] gzdLLzilambda11777R99;
  logic [0:0] callResR199;
  logic [106:0] gzdLLzilambda11786;
  logic [0:0] callResR200;
  logic [106:0] gzdLLzilambda11786R1;
  logic [0:0] callResR201;
  logic [106:0] gzdLLzilambda11786R2;
  logic [0:0] callResR202;
  logic [106:0] gzdLLzilambda11786R3;
  logic [0:0] callResR203;
  logic [106:0] gzdLLzilambda11786R4;
  logic [0:0] callResR204;
  logic [106:0] gzdLLzilambda11786R5;
  logic [0:0] callResR205;
  logic [106:0] gzdLLzilambda11786R6;
  logic [0:0] callResR206;
  logic [106:0] gzdLLzilambda11786R7;
  logic [0:0] callResR207;
  logic [106:0] gzdLLzilambda11786R8;
  logic [0:0] callResR208;
  logic [106:0] gzdLLzilambda11786R9;
  logic [0:0] callResR209;
  logic [106:0] gzdLLzilambda11786R10;
  logic [0:0] callResR210;
  logic [106:0] gzdLLzilambda11786R11;
  logic [0:0] callResR211;
  logic [106:0] gzdLLzilambda11786R12;
  logic [0:0] callResR212;
  logic [106:0] gzdLLzilambda11786R13;
  logic [0:0] callResR213;
  logic [106:0] gzdLLzilambda11786R14;
  logic [0:0] callResR214;
  logic [106:0] gzdLLzilambda11786R15;
  logic [0:0] callResR215;
  logic [106:0] gzdLLzilambda11786R16;
  logic [0:0] callResR216;
  logic [106:0] gzdLLzilambda11786R17;
  logic [0:0] callResR217;
  logic [106:0] gzdLLzilambda11786R18;
  logic [0:0] callResR218;
  logic [106:0] gzdLLzilambda11786R19;
  logic [0:0] callResR219;
  logic [106:0] gzdLLzilambda11786R20;
  logic [0:0] callResR220;
  logic [106:0] gzdLLzilambda11786R21;
  logic [0:0] callResR221;
  logic [106:0] gzdLLzilambda11786R22;
  logic [0:0] callResR222;
  logic [106:0] gzdLLzilambda11786R23;
  logic [0:0] callResR223;
  logic [106:0] gzdLLzilambda11786R24;
  logic [0:0] callResR224;
  logic [106:0] gzdLLzilambda11786R25;
  logic [0:0] callResR225;
  logic [106:0] gzdLLzilambda11786R26;
  logic [0:0] callResR226;
  logic [106:0] gzdLLzilambda11786R27;
  logic [0:0] callResR227;
  logic [106:0] gzdLLzilambda11786R28;
  logic [0:0] callResR228;
  logic [106:0] gzdLLzilambda11786R29;
  logic [0:0] callResR229;
  logic [106:0] gzdLLzilambda11786R30;
  logic [0:0] callResR230;
  logic [106:0] gzdLLzilambda11786R31;
  logic [0:0] callResR231;
  logic [106:0] gzdLLzilambda11786R32;
  logic [0:0] callResR232;
  logic [106:0] gzdLLzilambda11786R33;
  logic [0:0] callResR233;
  logic [106:0] gzdLLzilambda11786R34;
  logic [0:0] callResR234;
  logic [106:0] gzdLLzilambda11786R35;
  logic [0:0] callResR235;
  logic [106:0] gzdLLzilambda11786R36;
  logic [0:0] callResR236;
  logic [106:0] gzdLLzilambda11786R37;
  logic [0:0] callResR237;
  logic [106:0] gzdLLzilambda11786R38;
  logic [0:0] callResR238;
  logic [106:0] gzdLLzilambda11786R39;
  logic [0:0] callResR239;
  logic [106:0] gzdLLzilambda11786R40;
  logic [0:0] callResR240;
  logic [106:0] gzdLLzilambda11786R41;
  logic [0:0] callResR241;
  logic [106:0] gzdLLzilambda11786R42;
  logic [0:0] callResR242;
  logic [106:0] gzdLLzilambda11786R43;
  logic [0:0] callResR243;
  logic [106:0] gzdLLzilambda11786R44;
  logic [0:0] callResR244;
  logic [106:0] gzdLLzilambda11786R45;
  logic [0:0] callResR245;
  logic [106:0] gzdLLzilambda11786R46;
  logic [0:0] callResR246;
  logic [106:0] gzdLLzilambda11786R47;
  logic [0:0] callResR247;
  logic [106:0] gzdLLzilambda11786R48;
  logic [0:0] callResR248;
  logic [106:0] gzdLLzilambda11786R49;
  logic [0:0] callResR249;
  logic [106:0] gzdLLzilambda11786R50;
  logic [0:0] callResR250;
  logic [106:0] gzdLLzilambda11786R51;
  logic [0:0] callResR251;
  logic [106:0] gzdLLzilambda11786R52;
  logic [0:0] callResR252;
  logic [106:0] gzdLLzilambda11786R53;
  logic [0:0] callResR253;
  logic [106:0] gzdLLzilambda11786R54;
  logic [0:0] callResR254;
  logic [106:0] gzdLLzilambda11786R55;
  logic [0:0] callResR255;
  logic [106:0] gzdLLzilambda11786R56;
  logic [0:0] callResR256;
  logic [106:0] gzdLLzilambda11786R57;
  logic [0:0] callResR257;
  logic [106:0] gzdLLzilambda11786R58;
  logic [0:0] callResR258;
  logic [106:0] gzdLLzilambda11786R59;
  logic [0:0] callResR259;
  logic [106:0] gzdLLzilambda11786R60;
  logic [0:0] callResR260;
  logic [106:0] gzdLLzilambda11786R61;
  logic [0:0] callResR261;
  logic [106:0] gzdLLzilambda11786R62;
  logic [0:0] callResR262;
  logic [106:0] gzdLLzilambda11786R63;
  logic [0:0] callResR263;
  logic [106:0] gzdLLzilambda11786R64;
  logic [0:0] callResR264;
  logic [106:0] gzdLLzilambda11786R65;
  logic [0:0] callResR265;
  logic [106:0] gzdLLzilambda11786R66;
  logic [0:0] callResR266;
  logic [106:0] gzdLLzilambda11786R67;
  logic [0:0] callResR267;
  logic [106:0] gzdLLzilambda11786R68;
  logic [0:0] callResR268;
  logic [106:0] gzdLLzilambda11786R69;
  logic [0:0] callResR269;
  logic [106:0] gzdLLzilambda11786R70;
  logic [0:0] callResR270;
  logic [106:0] gzdLLzilambda11786R71;
  logic [0:0] callResR271;
  logic [106:0] gzdLLzilambda11786R72;
  logic [0:0] callResR272;
  logic [106:0] gzdLLzilambda11786R73;
  logic [0:0] callResR273;
  logic [106:0] gzdLLzilambda11786R74;
  logic [0:0] callResR274;
  logic [106:0] gzdLLzilambda11786R75;
  logic [0:0] callResR275;
  logic [106:0] gzdLLzilambda11786R76;
  logic [0:0] callResR276;
  logic [106:0] gzdLLzilambda11786R77;
  logic [0:0] callResR277;
  logic [106:0] gzdLLzilambda11786R78;
  logic [0:0] callResR278;
  logic [106:0] gzdLLzilambda11786R79;
  logic [0:0] callResR279;
  logic [106:0] gzdLLzilambda11786R80;
  logic [0:0] callResR280;
  logic [106:0] gzdLLzilambda11786R81;
  logic [0:0] callResR281;
  logic [106:0] gzdLLzilambda11786R82;
  logic [0:0] callResR282;
  logic [106:0] gzdLLzilambda11786R83;
  logic [0:0] callResR283;
  logic [106:0] gzdLLzilambda11786R84;
  logic [0:0] callResR284;
  logic [106:0] gzdLLzilambda11786R85;
  logic [0:0] callResR285;
  logic [106:0] gzdLLzilambda11786R86;
  logic [0:0] callResR286;
  logic [106:0] gzdLLzilambda11786R87;
  logic [0:0] callResR287;
  logic [106:0] gzdLLzilambda11786R88;
  logic [0:0] callResR288;
  logic [106:0] gzdLLzilambda11786R89;
  logic [0:0] callResR289;
  logic [106:0] gzdLLzilambda11786R90;
  logic [0:0] callResR290;
  logic [106:0] gzdLLzilambda11786R91;
  logic [0:0] callResR291;
  logic [106:0] gzdLLzilambda11786R92;
  logic [0:0] callResR292;
  logic [106:0] gzdLLzilambda11786R93;
  logic [0:0] callResR293;
  logic [106:0] gzdLLzilambda11786R94;
  logic [0:0] callResR294;
  logic [106:0] gzdLLzilambda11786R95;
  logic [0:0] callResR295;
  logic [106:0] gzdLLzilambda11786R96;
  logic [0:0] callResR296;
  logic [106:0] gzdLLzilambda11786R97;
  logic [0:0] callResR297;
  logic [106:0] gzdLLzilambda11786R98;
  logic [0:0] callResR298;
  logic [106:0] gzdLLzilambda11786R99;
  logic [0:0] callResR299;
  logic [106:0] gzdLLzilambda11795;
  logic [0:0] callResR300;
  logic [106:0] gzdLLzilambda11795R1;
  logic [0:0] callResR301;
  logic [106:0] gzdLLzilambda11795R2;
  logic [0:0] callResR302;
  logic [106:0] gzdLLzilambda11795R3;
  logic [0:0] callResR303;
  logic [106:0] gzdLLzilambda11795R4;
  logic [0:0] callResR304;
  logic [106:0] gzdLLzilambda11795R5;
  logic [0:0] callResR305;
  logic [106:0] gzdLLzilambda11795R6;
  logic [0:0] callResR306;
  logic [106:0] gzdLLzilambda11795R7;
  logic [0:0] callResR307;
  logic [106:0] gzdLLzilambda11795R8;
  logic [0:0] callResR308;
  logic [106:0] gzdLLzilambda11795R9;
  logic [0:0] callResR309;
  logic [106:0] gzdLLzilambda11795R10;
  logic [0:0] callResR310;
  logic [106:0] gzdLLzilambda11795R11;
  logic [0:0] callResR311;
  logic [106:0] gzdLLzilambda11795R12;
  logic [0:0] callResR312;
  logic [106:0] gzdLLzilambda11795R13;
  logic [0:0] callResR313;
  logic [106:0] gzdLLzilambda11795R14;
  logic [0:0] callResR314;
  logic [106:0] gzdLLzilambda11795R15;
  logic [0:0] callResR315;
  logic [106:0] gzdLLzilambda11795R16;
  logic [0:0] callResR316;
  logic [106:0] gzdLLzilambda11795R17;
  logic [0:0] callResR317;
  logic [106:0] gzdLLzilambda11795R18;
  logic [0:0] callResR318;
  logic [106:0] gzdLLzilambda11795R19;
  logic [0:0] callResR319;
  logic [106:0] gzdLLzilambda11795R20;
  logic [0:0] callResR320;
  logic [106:0] gzdLLzilambda11795R21;
  logic [0:0] callResR321;
  logic [106:0] gzdLLzilambda11795R22;
  logic [0:0] callResR322;
  logic [106:0] gzdLLzilambda11795R23;
  logic [0:0] callResR323;
  logic [106:0] gzdLLzilambda11795R24;
  logic [0:0] callResR324;
  logic [106:0] gzdLLzilambda11795R25;
  logic [0:0] callResR325;
  logic [106:0] gzdLLzilambda11795R26;
  logic [0:0] callResR326;
  logic [106:0] gzdLLzilambda11795R27;
  logic [0:0] callResR327;
  logic [106:0] gzdLLzilambda11795R28;
  logic [0:0] callResR328;
  logic [106:0] gzdLLzilambda11795R29;
  logic [0:0] callResR329;
  logic [106:0] gzdLLzilambda11795R30;
  logic [0:0] callResR330;
  logic [106:0] gzdLLzilambda11795R31;
  logic [0:0] callResR331;
  logic [106:0] gzdLLzilambda11795R32;
  logic [0:0] callResR332;
  logic [106:0] gzdLLzilambda11795R33;
  logic [0:0] callResR333;
  logic [106:0] gzdLLzilambda11795R34;
  logic [0:0] callResR334;
  logic [106:0] gzdLLzilambda11795R35;
  logic [0:0] callResR335;
  logic [106:0] gzdLLzilambda11795R36;
  logic [0:0] callResR336;
  logic [106:0] gzdLLzilambda11795R37;
  logic [0:0] callResR337;
  logic [106:0] gzdLLzilambda11795R38;
  logic [0:0] callResR338;
  logic [106:0] gzdLLzilambda11795R39;
  logic [0:0] callResR339;
  logic [106:0] gzdLLzilambda11795R40;
  logic [0:0] callResR340;
  logic [106:0] gzdLLzilambda11795R41;
  logic [0:0] callResR341;
  logic [106:0] gzdLLzilambda11795R42;
  logic [0:0] callResR342;
  logic [106:0] gzdLLzilambda11795R43;
  logic [0:0] callResR343;
  logic [106:0] gzdLLzilambda11795R44;
  logic [0:0] callResR344;
  logic [106:0] gzdLLzilambda11795R45;
  logic [0:0] callResR345;
  logic [106:0] gzdLLzilambda11795R46;
  logic [0:0] callResR346;
  logic [106:0] gzdLLzilambda11795R47;
  logic [0:0] callResR347;
  logic [106:0] gzdLLzilambda11795R48;
  logic [0:0] callResR348;
  logic [106:0] gzdLLzilambda11795R49;
  logic [0:0] callResR349;
  logic [106:0] gzdLLzilambda11795R50;
  logic [0:0] callResR350;
  logic [106:0] gzdLLzilambda11795R51;
  logic [0:0] callResR351;
  logic [106:0] gzdLLzilambda11795R52;
  logic [0:0] callResR352;
  logic [106:0] gzdLLzilambda11795R53;
  logic [0:0] callResR353;
  logic [106:0] gzdLLzilambda11795R54;
  logic [0:0] callResR354;
  logic [106:0] gzdLLzilambda11795R55;
  logic [0:0] callResR355;
  logic [106:0] gzdLLzilambda11795R56;
  logic [0:0] callResR356;
  logic [106:0] gzdLLzilambda11795R57;
  logic [0:0] callResR357;
  logic [106:0] gzdLLzilambda11795R58;
  logic [0:0] callResR358;
  logic [106:0] gzdLLzilambda11795R59;
  logic [0:0] callResR359;
  logic [106:0] gzdLLzilambda11795R60;
  logic [0:0] callResR360;
  logic [106:0] gzdLLzilambda11795R61;
  logic [0:0] callResR361;
  logic [106:0] gzdLLzilambda11795R62;
  logic [0:0] callResR362;
  logic [106:0] gzdLLzilambda11795R63;
  logic [0:0] callResR363;
  logic [106:0] gzdLLzilambda11795R64;
  logic [0:0] callResR364;
  logic [106:0] gzdLLzilambda11795R65;
  logic [0:0] callResR365;
  logic [106:0] gzdLLzilambda11795R66;
  logic [0:0] callResR366;
  logic [106:0] gzdLLzilambda11795R67;
  logic [0:0] callResR367;
  logic [106:0] gzdLLzilambda11795R68;
  logic [0:0] callResR368;
  logic [106:0] gzdLLzilambda11795R69;
  logic [0:0] callResR369;
  logic [106:0] gzdLLzilambda11795R70;
  logic [0:0] callResR370;
  logic [106:0] gzdLLzilambda11795R71;
  logic [0:0] callResR371;
  logic [106:0] gzdLLzilambda11795R72;
  logic [0:0] callResR372;
  logic [106:0] gzdLLzilambda11795R73;
  logic [0:0] callResR373;
  logic [106:0] gzdLLzilambda11795R74;
  logic [0:0] callResR374;
  logic [106:0] gzdLLzilambda11795R75;
  logic [0:0] callResR375;
  logic [106:0] gzdLLzilambda11795R76;
  logic [0:0] callResR376;
  logic [106:0] gzdLLzilambda11795R77;
  logic [0:0] callResR377;
  logic [106:0] gzdLLzilambda11795R78;
  logic [0:0] callResR378;
  logic [106:0] gzdLLzilambda11795R79;
  logic [0:0] callResR379;
  logic [106:0] gzdLLzilambda11795R80;
  logic [0:0] callResR380;
  logic [106:0] gzdLLzilambda11795R81;
  logic [0:0] callResR381;
  logic [106:0] gzdLLzilambda11795R82;
  logic [0:0] callResR382;
  logic [106:0] gzdLLzilambda11795R83;
  logic [0:0] callResR383;
  logic [106:0] gzdLLzilambda11795R84;
  logic [0:0] callResR384;
  logic [106:0] gzdLLzilambda11795R85;
  logic [0:0] callResR385;
  logic [106:0] gzdLLzilambda11795R86;
  logic [0:0] callResR386;
  logic [106:0] gzdLLzilambda11795R87;
  logic [0:0] callResR387;
  logic [106:0] gzdLLzilambda11795R88;
  logic [0:0] callResR388;
  logic [106:0] gzdLLzilambda11795R89;
  logic [0:0] callResR389;
  logic [106:0] gzdLLzilambda11795R90;
  logic [0:0] callResR390;
  logic [106:0] gzdLLzilambda11795R91;
  logic [0:0] callResR391;
  logic [106:0] gzdLLzilambda11795R92;
  logic [0:0] callResR392;
  logic [106:0] gzdLLzilambda11795R93;
  logic [0:0] callResR393;
  logic [106:0] gzdLLzilambda11795R94;
  logic [0:0] callResR394;
  logic [106:0] gzdLLzilambda11795R95;
  logic [0:0] callResR395;
  logic [106:0] gzdLLzilambda11795R96;
  logic [0:0] callResR396;
  logic [106:0] gzdLLzilambda11795R97;
  logic [0:0] callResR397;
  logic [106:0] gzdLLzilambda11795R98;
  logic [0:0] callResR398;
  logic [106:0] gzdLLzilambda11795R99;
  logic [0:0] callResR399;
  assign gMainzidev = arg0;
  assign gzdLLzilambda11768 = {gMainzidev[99:0], 7'h00};
  zdLLzilambda11768  zdLLzilambda11768 (gzdLLzilambda11768[106:7], gzdLLzilambda11768[6:0], callRes);
  assign gzdLLzilambda11768R1 = {gMainzidev[99:0], 7'h01};
  zdLLzilambda11768  zdLLzilambda11768R1 (gzdLLzilambda11768R1[106:7], gzdLLzilambda11768R1[6:0], callResR1);
  assign gzdLLzilambda11768R2 = {gMainzidev[99:0], 7'h02};
  zdLLzilambda11768  zdLLzilambda11768R2 (gzdLLzilambda11768R2[106:7], gzdLLzilambda11768R2[6:0], callResR2);
  assign gzdLLzilambda11768R3 = {gMainzidev[99:0], 7'h03};
  zdLLzilambda11768  zdLLzilambda11768R3 (gzdLLzilambda11768R3[106:7], gzdLLzilambda11768R3[6:0], callResR3);
  assign gzdLLzilambda11768R4 = {gMainzidev[99:0], 7'h04};
  zdLLzilambda11768  zdLLzilambda11768R4 (gzdLLzilambda11768R4[106:7], gzdLLzilambda11768R4[6:0], callResR4);
  assign gzdLLzilambda11768R5 = {gMainzidev[99:0], 7'h05};
  zdLLzilambda11768  zdLLzilambda11768R5 (gzdLLzilambda11768R5[106:7], gzdLLzilambda11768R5[6:0], callResR5);
  assign gzdLLzilambda11768R6 = {gMainzidev[99:0], 7'h06};
  zdLLzilambda11768  zdLLzilambda11768R6 (gzdLLzilambda11768R6[106:7], gzdLLzilambda11768R6[6:0], callResR6);
  assign gzdLLzilambda11768R7 = {gMainzidev[99:0], 7'h07};
  zdLLzilambda11768  zdLLzilambda11768R7 (gzdLLzilambda11768R7[106:7], gzdLLzilambda11768R7[6:0], callResR7);
  assign gzdLLzilambda11768R8 = {gMainzidev[99:0], 7'h08};
  zdLLzilambda11768  zdLLzilambda11768R8 (gzdLLzilambda11768R8[106:7], gzdLLzilambda11768R8[6:0], callResR8);
  assign gzdLLzilambda11768R9 = {gMainzidev[99:0], 7'h09};
  zdLLzilambda11768  zdLLzilambda11768R9 (gzdLLzilambda11768R9[106:7], gzdLLzilambda11768R9[6:0], callResR9);
  assign gzdLLzilambda11768R10 = {gMainzidev[99:0], 7'h0a};
  zdLLzilambda11768  zdLLzilambda11768R10 (gzdLLzilambda11768R10[106:7], gzdLLzilambda11768R10[6:0], callResR10);
  assign gzdLLzilambda11768R11 = {gMainzidev[99:0], 7'h0b};
  zdLLzilambda11768  zdLLzilambda11768R11 (gzdLLzilambda11768R11[106:7], gzdLLzilambda11768R11[6:0], callResR11);
  assign gzdLLzilambda11768R12 = {gMainzidev[99:0], 7'h0c};
  zdLLzilambda11768  zdLLzilambda11768R12 (gzdLLzilambda11768R12[106:7], gzdLLzilambda11768R12[6:0], callResR12);
  assign gzdLLzilambda11768R13 = {gMainzidev[99:0], 7'h0d};
  zdLLzilambda11768  zdLLzilambda11768R13 (gzdLLzilambda11768R13[106:7], gzdLLzilambda11768R13[6:0], callResR13);
  assign gzdLLzilambda11768R14 = {gMainzidev[99:0], 7'h0e};
  zdLLzilambda11768  zdLLzilambda11768R14 (gzdLLzilambda11768R14[106:7], gzdLLzilambda11768R14[6:0], callResR14);
  assign gzdLLzilambda11768R15 = {gMainzidev[99:0], 7'h0f};
  zdLLzilambda11768  zdLLzilambda11768R15 (gzdLLzilambda11768R15[106:7], gzdLLzilambda11768R15[6:0], callResR15);
  assign gzdLLzilambda11768R16 = {gMainzidev[99:0], 7'h10};
  zdLLzilambda11768  zdLLzilambda11768R16 (gzdLLzilambda11768R16[106:7], gzdLLzilambda11768R16[6:0], callResR16);
  assign gzdLLzilambda11768R17 = {gMainzidev[99:0], 7'h11};
  zdLLzilambda11768  zdLLzilambda11768R17 (gzdLLzilambda11768R17[106:7], gzdLLzilambda11768R17[6:0], callResR17);
  assign gzdLLzilambda11768R18 = {gMainzidev[99:0], 7'h12};
  zdLLzilambda11768  zdLLzilambda11768R18 (gzdLLzilambda11768R18[106:7], gzdLLzilambda11768R18[6:0], callResR18);
  assign gzdLLzilambda11768R19 = {gMainzidev[99:0], 7'h13};
  zdLLzilambda11768  zdLLzilambda11768R19 (gzdLLzilambda11768R19[106:7], gzdLLzilambda11768R19[6:0], callResR19);
  assign gzdLLzilambda11768R20 = {gMainzidev[99:0], 7'h14};
  zdLLzilambda11768  zdLLzilambda11768R20 (gzdLLzilambda11768R20[106:7], gzdLLzilambda11768R20[6:0], callResR20);
  assign gzdLLzilambda11768R21 = {gMainzidev[99:0], 7'h15};
  zdLLzilambda11768  zdLLzilambda11768R21 (gzdLLzilambda11768R21[106:7], gzdLLzilambda11768R21[6:0], callResR21);
  assign gzdLLzilambda11768R22 = {gMainzidev[99:0], 7'h16};
  zdLLzilambda11768  zdLLzilambda11768R22 (gzdLLzilambda11768R22[106:7], gzdLLzilambda11768R22[6:0], callResR22);
  assign gzdLLzilambda11768R23 = {gMainzidev[99:0], 7'h17};
  zdLLzilambda11768  zdLLzilambda11768R23 (gzdLLzilambda11768R23[106:7], gzdLLzilambda11768R23[6:0], callResR23);
  assign gzdLLzilambda11768R24 = {gMainzidev[99:0], 7'h18};
  zdLLzilambda11768  zdLLzilambda11768R24 (gzdLLzilambda11768R24[106:7], gzdLLzilambda11768R24[6:0], callResR24);
  assign gzdLLzilambda11768R25 = {gMainzidev[99:0], 7'h19};
  zdLLzilambda11768  zdLLzilambda11768R25 (gzdLLzilambda11768R25[106:7], gzdLLzilambda11768R25[6:0], callResR25);
  assign gzdLLzilambda11768R26 = {gMainzidev[99:0], 7'h1a};
  zdLLzilambda11768  zdLLzilambda11768R26 (gzdLLzilambda11768R26[106:7], gzdLLzilambda11768R26[6:0], callResR26);
  assign gzdLLzilambda11768R27 = {gMainzidev[99:0], 7'h1b};
  zdLLzilambda11768  zdLLzilambda11768R27 (gzdLLzilambda11768R27[106:7], gzdLLzilambda11768R27[6:0], callResR27);
  assign gzdLLzilambda11768R28 = {gMainzidev[99:0], 7'h1c};
  zdLLzilambda11768  zdLLzilambda11768R28 (gzdLLzilambda11768R28[106:7], gzdLLzilambda11768R28[6:0], callResR28);
  assign gzdLLzilambda11768R29 = {gMainzidev[99:0], 7'h1d};
  zdLLzilambda11768  zdLLzilambda11768R29 (gzdLLzilambda11768R29[106:7], gzdLLzilambda11768R29[6:0], callResR29);
  assign gzdLLzilambda11768R30 = {gMainzidev[99:0], 7'h1e};
  zdLLzilambda11768  zdLLzilambda11768R30 (gzdLLzilambda11768R30[106:7], gzdLLzilambda11768R30[6:0], callResR30);
  assign gzdLLzilambda11768R31 = {gMainzidev[99:0], 7'h1f};
  zdLLzilambda11768  zdLLzilambda11768R31 (gzdLLzilambda11768R31[106:7], gzdLLzilambda11768R31[6:0], callResR31);
  assign gzdLLzilambda11768R32 = {gMainzidev[99:0], 7'h20};
  zdLLzilambda11768  zdLLzilambda11768R32 (gzdLLzilambda11768R32[106:7], gzdLLzilambda11768R32[6:0], callResR32);
  assign gzdLLzilambda11768R33 = {gMainzidev[99:0], 7'h21};
  zdLLzilambda11768  zdLLzilambda11768R33 (gzdLLzilambda11768R33[106:7], gzdLLzilambda11768R33[6:0], callResR33);
  assign gzdLLzilambda11768R34 = {gMainzidev[99:0], 7'h22};
  zdLLzilambda11768  zdLLzilambda11768R34 (gzdLLzilambda11768R34[106:7], gzdLLzilambda11768R34[6:0], callResR34);
  assign gzdLLzilambda11768R35 = {gMainzidev[99:0], 7'h23};
  zdLLzilambda11768  zdLLzilambda11768R35 (gzdLLzilambda11768R35[106:7], gzdLLzilambda11768R35[6:0], callResR35);
  assign gzdLLzilambda11768R36 = {gMainzidev[99:0], 7'h24};
  zdLLzilambda11768  zdLLzilambda11768R36 (gzdLLzilambda11768R36[106:7], gzdLLzilambda11768R36[6:0], callResR36);
  assign gzdLLzilambda11768R37 = {gMainzidev[99:0], 7'h25};
  zdLLzilambda11768  zdLLzilambda11768R37 (gzdLLzilambda11768R37[106:7], gzdLLzilambda11768R37[6:0], callResR37);
  assign gzdLLzilambda11768R38 = {gMainzidev[99:0], 7'h26};
  zdLLzilambda11768  zdLLzilambda11768R38 (gzdLLzilambda11768R38[106:7], gzdLLzilambda11768R38[6:0], callResR38);
  assign gzdLLzilambda11768R39 = {gMainzidev[99:0], 7'h27};
  zdLLzilambda11768  zdLLzilambda11768R39 (gzdLLzilambda11768R39[106:7], gzdLLzilambda11768R39[6:0], callResR39);
  assign gzdLLzilambda11768R40 = {gMainzidev[99:0], 7'h28};
  zdLLzilambda11768  zdLLzilambda11768R40 (gzdLLzilambda11768R40[106:7], gzdLLzilambda11768R40[6:0], callResR40);
  assign gzdLLzilambda11768R41 = {gMainzidev[99:0], 7'h29};
  zdLLzilambda11768  zdLLzilambda11768R41 (gzdLLzilambda11768R41[106:7], gzdLLzilambda11768R41[6:0], callResR41);
  assign gzdLLzilambda11768R42 = {gMainzidev[99:0], 7'h2a};
  zdLLzilambda11768  zdLLzilambda11768R42 (gzdLLzilambda11768R42[106:7], gzdLLzilambda11768R42[6:0], callResR42);
  assign gzdLLzilambda11768R43 = {gMainzidev[99:0], 7'h2b};
  zdLLzilambda11768  zdLLzilambda11768R43 (gzdLLzilambda11768R43[106:7], gzdLLzilambda11768R43[6:0], callResR43);
  assign gzdLLzilambda11768R44 = {gMainzidev[99:0], 7'h2c};
  zdLLzilambda11768  zdLLzilambda11768R44 (gzdLLzilambda11768R44[106:7], gzdLLzilambda11768R44[6:0], callResR44);
  assign gzdLLzilambda11768R45 = {gMainzidev[99:0], 7'h2d};
  zdLLzilambda11768  zdLLzilambda11768R45 (gzdLLzilambda11768R45[106:7], gzdLLzilambda11768R45[6:0], callResR45);
  assign gzdLLzilambda11768R46 = {gMainzidev[99:0], 7'h2e};
  zdLLzilambda11768  zdLLzilambda11768R46 (gzdLLzilambda11768R46[106:7], gzdLLzilambda11768R46[6:0], callResR46);
  assign gzdLLzilambda11768R47 = {gMainzidev[99:0], 7'h2f};
  zdLLzilambda11768  zdLLzilambda11768R47 (gzdLLzilambda11768R47[106:7], gzdLLzilambda11768R47[6:0], callResR47);
  assign gzdLLzilambda11768R48 = {gMainzidev[99:0], 7'h30};
  zdLLzilambda11768  zdLLzilambda11768R48 (gzdLLzilambda11768R48[106:7], gzdLLzilambda11768R48[6:0], callResR48);
  assign gzdLLzilambda11768R49 = {gMainzidev[99:0], 7'h31};
  zdLLzilambda11768  zdLLzilambda11768R49 (gzdLLzilambda11768R49[106:7], gzdLLzilambda11768R49[6:0], callResR49);
  assign gzdLLzilambda11768R50 = {gMainzidev[99:0], 7'h32};
  zdLLzilambda11768  zdLLzilambda11768R50 (gzdLLzilambda11768R50[106:7], gzdLLzilambda11768R50[6:0], callResR50);
  assign gzdLLzilambda11768R51 = {gMainzidev[99:0], 7'h33};
  zdLLzilambda11768  zdLLzilambda11768R51 (gzdLLzilambda11768R51[106:7], gzdLLzilambda11768R51[6:0], callResR51);
  assign gzdLLzilambda11768R52 = {gMainzidev[99:0], 7'h34};
  zdLLzilambda11768  zdLLzilambda11768R52 (gzdLLzilambda11768R52[106:7], gzdLLzilambda11768R52[6:0], callResR52);
  assign gzdLLzilambda11768R53 = {gMainzidev[99:0], 7'h35};
  zdLLzilambda11768  zdLLzilambda11768R53 (gzdLLzilambda11768R53[106:7], gzdLLzilambda11768R53[6:0], callResR53);
  assign gzdLLzilambda11768R54 = {gMainzidev[99:0], 7'h36};
  zdLLzilambda11768  zdLLzilambda11768R54 (gzdLLzilambda11768R54[106:7], gzdLLzilambda11768R54[6:0], callResR54);
  assign gzdLLzilambda11768R55 = {gMainzidev[99:0], 7'h37};
  zdLLzilambda11768  zdLLzilambda11768R55 (gzdLLzilambda11768R55[106:7], gzdLLzilambda11768R55[6:0], callResR55);
  assign gzdLLzilambda11768R56 = {gMainzidev[99:0], 7'h38};
  zdLLzilambda11768  zdLLzilambda11768R56 (gzdLLzilambda11768R56[106:7], gzdLLzilambda11768R56[6:0], callResR56);
  assign gzdLLzilambda11768R57 = {gMainzidev[99:0], 7'h39};
  zdLLzilambda11768  zdLLzilambda11768R57 (gzdLLzilambda11768R57[106:7], gzdLLzilambda11768R57[6:0], callResR57);
  assign gzdLLzilambda11768R58 = {gMainzidev[99:0], 7'h3a};
  zdLLzilambda11768  zdLLzilambda11768R58 (gzdLLzilambda11768R58[106:7], gzdLLzilambda11768R58[6:0], callResR58);
  assign gzdLLzilambda11768R59 = {gMainzidev[99:0], 7'h3b};
  zdLLzilambda11768  zdLLzilambda11768R59 (gzdLLzilambda11768R59[106:7], gzdLLzilambda11768R59[6:0], callResR59);
  assign gzdLLzilambda11768R60 = {gMainzidev[99:0], 7'h3c};
  zdLLzilambda11768  zdLLzilambda11768R60 (gzdLLzilambda11768R60[106:7], gzdLLzilambda11768R60[6:0], callResR60);
  assign gzdLLzilambda11768R61 = {gMainzidev[99:0], 7'h3d};
  zdLLzilambda11768  zdLLzilambda11768R61 (gzdLLzilambda11768R61[106:7], gzdLLzilambda11768R61[6:0], callResR61);
  assign gzdLLzilambda11768R62 = {gMainzidev[99:0], 7'h3e};
  zdLLzilambda11768  zdLLzilambda11768R62 (gzdLLzilambda11768R62[106:7], gzdLLzilambda11768R62[6:0], callResR62);
  assign gzdLLzilambda11768R63 = {gMainzidev[99:0], 7'h3f};
  zdLLzilambda11768  zdLLzilambda11768R63 (gzdLLzilambda11768R63[106:7], gzdLLzilambda11768R63[6:0], callResR63);
  assign gzdLLzilambda11768R64 = {gMainzidev[99:0], 7'h40};
  zdLLzilambda11768  zdLLzilambda11768R64 (gzdLLzilambda11768R64[106:7], gzdLLzilambda11768R64[6:0], callResR64);
  assign gzdLLzilambda11768R65 = {gMainzidev[99:0], 7'h41};
  zdLLzilambda11768  zdLLzilambda11768R65 (gzdLLzilambda11768R65[106:7], gzdLLzilambda11768R65[6:0], callResR65);
  assign gzdLLzilambda11768R66 = {gMainzidev[99:0], 7'h42};
  zdLLzilambda11768  zdLLzilambda11768R66 (gzdLLzilambda11768R66[106:7], gzdLLzilambda11768R66[6:0], callResR66);
  assign gzdLLzilambda11768R67 = {gMainzidev[99:0], 7'h43};
  zdLLzilambda11768  zdLLzilambda11768R67 (gzdLLzilambda11768R67[106:7], gzdLLzilambda11768R67[6:0], callResR67);
  assign gzdLLzilambda11768R68 = {gMainzidev[99:0], 7'h44};
  zdLLzilambda11768  zdLLzilambda11768R68 (gzdLLzilambda11768R68[106:7], gzdLLzilambda11768R68[6:0], callResR68);
  assign gzdLLzilambda11768R69 = {gMainzidev[99:0], 7'h45};
  zdLLzilambda11768  zdLLzilambda11768R69 (gzdLLzilambda11768R69[106:7], gzdLLzilambda11768R69[6:0], callResR69);
  assign gzdLLzilambda11768R70 = {gMainzidev[99:0], 7'h46};
  zdLLzilambda11768  zdLLzilambda11768R70 (gzdLLzilambda11768R70[106:7], gzdLLzilambda11768R70[6:0], callResR70);
  assign gzdLLzilambda11768R71 = {gMainzidev[99:0], 7'h47};
  zdLLzilambda11768  zdLLzilambda11768R71 (gzdLLzilambda11768R71[106:7], gzdLLzilambda11768R71[6:0], callResR71);
  assign gzdLLzilambda11768R72 = {gMainzidev[99:0], 7'h48};
  zdLLzilambda11768  zdLLzilambda11768R72 (gzdLLzilambda11768R72[106:7], gzdLLzilambda11768R72[6:0], callResR72);
  assign gzdLLzilambda11768R73 = {gMainzidev[99:0], 7'h49};
  zdLLzilambda11768  zdLLzilambda11768R73 (gzdLLzilambda11768R73[106:7], gzdLLzilambda11768R73[6:0], callResR73);
  assign gzdLLzilambda11768R74 = {gMainzidev[99:0], 7'h4a};
  zdLLzilambda11768  zdLLzilambda11768R74 (gzdLLzilambda11768R74[106:7], gzdLLzilambda11768R74[6:0], callResR74);
  assign gzdLLzilambda11768R75 = {gMainzidev[99:0], 7'h4b};
  zdLLzilambda11768  zdLLzilambda11768R75 (gzdLLzilambda11768R75[106:7], gzdLLzilambda11768R75[6:0], callResR75);
  assign gzdLLzilambda11768R76 = {gMainzidev[99:0], 7'h4c};
  zdLLzilambda11768  zdLLzilambda11768R76 (gzdLLzilambda11768R76[106:7], gzdLLzilambda11768R76[6:0], callResR76);
  assign gzdLLzilambda11768R77 = {gMainzidev[99:0], 7'h4d};
  zdLLzilambda11768  zdLLzilambda11768R77 (gzdLLzilambda11768R77[106:7], gzdLLzilambda11768R77[6:0], callResR77);
  assign gzdLLzilambda11768R78 = {gMainzidev[99:0], 7'h4e};
  zdLLzilambda11768  zdLLzilambda11768R78 (gzdLLzilambda11768R78[106:7], gzdLLzilambda11768R78[6:0], callResR78);
  assign gzdLLzilambda11768R79 = {gMainzidev[99:0], 7'h4f};
  zdLLzilambda11768  zdLLzilambda11768R79 (gzdLLzilambda11768R79[106:7], gzdLLzilambda11768R79[6:0], callResR79);
  assign gzdLLzilambda11768R80 = {gMainzidev[99:0], 7'h50};
  zdLLzilambda11768  zdLLzilambda11768R80 (gzdLLzilambda11768R80[106:7], gzdLLzilambda11768R80[6:0], callResR80);
  assign gzdLLzilambda11768R81 = {gMainzidev[99:0], 7'h51};
  zdLLzilambda11768  zdLLzilambda11768R81 (gzdLLzilambda11768R81[106:7], gzdLLzilambda11768R81[6:0], callResR81);
  assign gzdLLzilambda11768R82 = {gMainzidev[99:0], 7'h52};
  zdLLzilambda11768  zdLLzilambda11768R82 (gzdLLzilambda11768R82[106:7], gzdLLzilambda11768R82[6:0], callResR82);
  assign gzdLLzilambda11768R83 = {gMainzidev[99:0], 7'h53};
  zdLLzilambda11768  zdLLzilambda11768R83 (gzdLLzilambda11768R83[106:7], gzdLLzilambda11768R83[6:0], callResR83);
  assign gzdLLzilambda11768R84 = {gMainzidev[99:0], 7'h54};
  zdLLzilambda11768  zdLLzilambda11768R84 (gzdLLzilambda11768R84[106:7], gzdLLzilambda11768R84[6:0], callResR84);
  assign gzdLLzilambda11768R85 = {gMainzidev[99:0], 7'h55};
  zdLLzilambda11768  zdLLzilambda11768R85 (gzdLLzilambda11768R85[106:7], gzdLLzilambda11768R85[6:0], callResR85);
  assign gzdLLzilambda11768R86 = {gMainzidev[99:0], 7'h56};
  zdLLzilambda11768  zdLLzilambda11768R86 (gzdLLzilambda11768R86[106:7], gzdLLzilambda11768R86[6:0], callResR86);
  assign gzdLLzilambda11768R87 = {gMainzidev[99:0], 7'h57};
  zdLLzilambda11768  zdLLzilambda11768R87 (gzdLLzilambda11768R87[106:7], gzdLLzilambda11768R87[6:0], callResR87);
  assign gzdLLzilambda11768R88 = {gMainzidev[99:0], 7'h58};
  zdLLzilambda11768  zdLLzilambda11768R88 (gzdLLzilambda11768R88[106:7], gzdLLzilambda11768R88[6:0], callResR88);
  assign gzdLLzilambda11768R89 = {gMainzidev[99:0], 7'h59};
  zdLLzilambda11768  zdLLzilambda11768R89 (gzdLLzilambda11768R89[106:7], gzdLLzilambda11768R89[6:0], callResR89);
  assign gzdLLzilambda11768R90 = {gMainzidev[99:0], 7'h5a};
  zdLLzilambda11768  zdLLzilambda11768R90 (gzdLLzilambda11768R90[106:7], gzdLLzilambda11768R90[6:0], callResR90);
  assign gzdLLzilambda11768R91 = {gMainzidev[99:0], 7'h5b};
  zdLLzilambda11768  zdLLzilambda11768R91 (gzdLLzilambda11768R91[106:7], gzdLLzilambda11768R91[6:0], callResR91);
  assign gzdLLzilambda11768R92 = {gMainzidev[99:0], 7'h5c};
  zdLLzilambda11768  zdLLzilambda11768R92 (gzdLLzilambda11768R92[106:7], gzdLLzilambda11768R92[6:0], callResR92);
  assign gzdLLzilambda11768R93 = {gMainzidev[99:0], 7'h5d};
  zdLLzilambda11768  zdLLzilambda11768R93 (gzdLLzilambda11768R93[106:7], gzdLLzilambda11768R93[6:0], callResR93);
  assign gzdLLzilambda11768R94 = {gMainzidev[99:0], 7'h5e};
  zdLLzilambda11768  zdLLzilambda11768R94 (gzdLLzilambda11768R94[106:7], gzdLLzilambda11768R94[6:0], callResR94);
  assign gzdLLzilambda11768R95 = {gMainzidev[99:0], 7'h5f};
  zdLLzilambda11768  zdLLzilambda11768R95 (gzdLLzilambda11768R95[106:7], gzdLLzilambda11768R95[6:0], callResR95);
  assign gzdLLzilambda11768R96 = {gMainzidev[99:0], 7'h60};
  zdLLzilambda11768  zdLLzilambda11768R96 (gzdLLzilambda11768R96[106:7], gzdLLzilambda11768R96[6:0], callResR96);
  assign gzdLLzilambda11768R97 = {gMainzidev[99:0], 7'h61};
  zdLLzilambda11768  zdLLzilambda11768R97 (gzdLLzilambda11768R97[106:7], gzdLLzilambda11768R97[6:0], callResR97);
  assign gzdLLzilambda11768R98 = {gMainzidev[99:0], 7'h62};
  zdLLzilambda11768  zdLLzilambda11768R98 (gzdLLzilambda11768R98[106:7], gzdLLzilambda11768R98[6:0], callResR98);
  assign gzdLLzilambda11768R99 = {gMainzidev[99:0], 7'h63};
  zdLLzilambda11768  zdLLzilambda11768R99 (gzdLLzilambda11768R99[106:7], gzdLLzilambda11768R99[6:0], callResR99);
  assign gzdLLzilambda11777 = {gMainzidev[99:0], 7'h00};
  zdLLzilambda11777  zdLLzilambda11777 (gzdLLzilambda11777[106:7], gzdLLzilambda11777[6:0], callResR100);
  assign gzdLLzilambda11777R1 = {gMainzidev[99:0], 7'h01};
  zdLLzilambda11777  zdLLzilambda11777R1 (gzdLLzilambda11777R1[106:7], gzdLLzilambda11777R1[6:0], callResR101);
  assign gzdLLzilambda11777R2 = {gMainzidev[99:0], 7'h02};
  zdLLzilambda11777  zdLLzilambda11777R2 (gzdLLzilambda11777R2[106:7], gzdLLzilambda11777R2[6:0], callResR102);
  assign gzdLLzilambda11777R3 = {gMainzidev[99:0], 7'h03};
  zdLLzilambda11777  zdLLzilambda11777R3 (gzdLLzilambda11777R3[106:7], gzdLLzilambda11777R3[6:0], callResR103);
  assign gzdLLzilambda11777R4 = {gMainzidev[99:0], 7'h04};
  zdLLzilambda11777  zdLLzilambda11777R4 (gzdLLzilambda11777R4[106:7], gzdLLzilambda11777R4[6:0], callResR104);
  assign gzdLLzilambda11777R5 = {gMainzidev[99:0], 7'h05};
  zdLLzilambda11777  zdLLzilambda11777R5 (gzdLLzilambda11777R5[106:7], gzdLLzilambda11777R5[6:0], callResR105);
  assign gzdLLzilambda11777R6 = {gMainzidev[99:0], 7'h06};
  zdLLzilambda11777  zdLLzilambda11777R6 (gzdLLzilambda11777R6[106:7], gzdLLzilambda11777R6[6:0], callResR106);
  assign gzdLLzilambda11777R7 = {gMainzidev[99:0], 7'h07};
  zdLLzilambda11777  zdLLzilambda11777R7 (gzdLLzilambda11777R7[106:7], gzdLLzilambda11777R7[6:0], callResR107);
  assign gzdLLzilambda11777R8 = {gMainzidev[99:0], 7'h08};
  zdLLzilambda11777  zdLLzilambda11777R8 (gzdLLzilambda11777R8[106:7], gzdLLzilambda11777R8[6:0], callResR108);
  assign gzdLLzilambda11777R9 = {gMainzidev[99:0], 7'h09};
  zdLLzilambda11777  zdLLzilambda11777R9 (gzdLLzilambda11777R9[106:7], gzdLLzilambda11777R9[6:0], callResR109);
  assign gzdLLzilambda11777R10 = {gMainzidev[99:0], 7'h0a};
  zdLLzilambda11777  zdLLzilambda11777R10 (gzdLLzilambda11777R10[106:7], gzdLLzilambda11777R10[6:0], callResR110);
  assign gzdLLzilambda11777R11 = {gMainzidev[99:0], 7'h0b};
  zdLLzilambda11777  zdLLzilambda11777R11 (gzdLLzilambda11777R11[106:7], gzdLLzilambda11777R11[6:0], callResR111);
  assign gzdLLzilambda11777R12 = {gMainzidev[99:0], 7'h0c};
  zdLLzilambda11777  zdLLzilambda11777R12 (gzdLLzilambda11777R12[106:7], gzdLLzilambda11777R12[6:0], callResR112);
  assign gzdLLzilambda11777R13 = {gMainzidev[99:0], 7'h0d};
  zdLLzilambda11777  zdLLzilambda11777R13 (gzdLLzilambda11777R13[106:7], gzdLLzilambda11777R13[6:0], callResR113);
  assign gzdLLzilambda11777R14 = {gMainzidev[99:0], 7'h0e};
  zdLLzilambda11777  zdLLzilambda11777R14 (gzdLLzilambda11777R14[106:7], gzdLLzilambda11777R14[6:0], callResR114);
  assign gzdLLzilambda11777R15 = {gMainzidev[99:0], 7'h0f};
  zdLLzilambda11777  zdLLzilambda11777R15 (gzdLLzilambda11777R15[106:7], gzdLLzilambda11777R15[6:0], callResR115);
  assign gzdLLzilambda11777R16 = {gMainzidev[99:0], 7'h10};
  zdLLzilambda11777  zdLLzilambda11777R16 (gzdLLzilambda11777R16[106:7], gzdLLzilambda11777R16[6:0], callResR116);
  assign gzdLLzilambda11777R17 = {gMainzidev[99:0], 7'h11};
  zdLLzilambda11777  zdLLzilambda11777R17 (gzdLLzilambda11777R17[106:7], gzdLLzilambda11777R17[6:0], callResR117);
  assign gzdLLzilambda11777R18 = {gMainzidev[99:0], 7'h12};
  zdLLzilambda11777  zdLLzilambda11777R18 (gzdLLzilambda11777R18[106:7], gzdLLzilambda11777R18[6:0], callResR118);
  assign gzdLLzilambda11777R19 = {gMainzidev[99:0], 7'h13};
  zdLLzilambda11777  zdLLzilambda11777R19 (gzdLLzilambda11777R19[106:7], gzdLLzilambda11777R19[6:0], callResR119);
  assign gzdLLzilambda11777R20 = {gMainzidev[99:0], 7'h14};
  zdLLzilambda11777  zdLLzilambda11777R20 (gzdLLzilambda11777R20[106:7], gzdLLzilambda11777R20[6:0], callResR120);
  assign gzdLLzilambda11777R21 = {gMainzidev[99:0], 7'h15};
  zdLLzilambda11777  zdLLzilambda11777R21 (gzdLLzilambda11777R21[106:7], gzdLLzilambda11777R21[6:0], callResR121);
  assign gzdLLzilambda11777R22 = {gMainzidev[99:0], 7'h16};
  zdLLzilambda11777  zdLLzilambda11777R22 (gzdLLzilambda11777R22[106:7], gzdLLzilambda11777R22[6:0], callResR122);
  assign gzdLLzilambda11777R23 = {gMainzidev[99:0], 7'h17};
  zdLLzilambda11777  zdLLzilambda11777R23 (gzdLLzilambda11777R23[106:7], gzdLLzilambda11777R23[6:0], callResR123);
  assign gzdLLzilambda11777R24 = {gMainzidev[99:0], 7'h18};
  zdLLzilambda11777  zdLLzilambda11777R24 (gzdLLzilambda11777R24[106:7], gzdLLzilambda11777R24[6:0], callResR124);
  assign gzdLLzilambda11777R25 = {gMainzidev[99:0], 7'h19};
  zdLLzilambda11777  zdLLzilambda11777R25 (gzdLLzilambda11777R25[106:7], gzdLLzilambda11777R25[6:0], callResR125);
  assign gzdLLzilambda11777R26 = {gMainzidev[99:0], 7'h1a};
  zdLLzilambda11777  zdLLzilambda11777R26 (gzdLLzilambda11777R26[106:7], gzdLLzilambda11777R26[6:0], callResR126);
  assign gzdLLzilambda11777R27 = {gMainzidev[99:0], 7'h1b};
  zdLLzilambda11777  zdLLzilambda11777R27 (gzdLLzilambda11777R27[106:7], gzdLLzilambda11777R27[6:0], callResR127);
  assign gzdLLzilambda11777R28 = {gMainzidev[99:0], 7'h1c};
  zdLLzilambda11777  zdLLzilambda11777R28 (gzdLLzilambda11777R28[106:7], gzdLLzilambda11777R28[6:0], callResR128);
  assign gzdLLzilambda11777R29 = {gMainzidev[99:0], 7'h1d};
  zdLLzilambda11777  zdLLzilambda11777R29 (gzdLLzilambda11777R29[106:7], gzdLLzilambda11777R29[6:0], callResR129);
  assign gzdLLzilambda11777R30 = {gMainzidev[99:0], 7'h1e};
  zdLLzilambda11777  zdLLzilambda11777R30 (gzdLLzilambda11777R30[106:7], gzdLLzilambda11777R30[6:0], callResR130);
  assign gzdLLzilambda11777R31 = {gMainzidev[99:0], 7'h1f};
  zdLLzilambda11777  zdLLzilambda11777R31 (gzdLLzilambda11777R31[106:7], gzdLLzilambda11777R31[6:0], callResR131);
  assign gzdLLzilambda11777R32 = {gMainzidev[99:0], 7'h20};
  zdLLzilambda11777  zdLLzilambda11777R32 (gzdLLzilambda11777R32[106:7], gzdLLzilambda11777R32[6:0], callResR132);
  assign gzdLLzilambda11777R33 = {gMainzidev[99:0], 7'h21};
  zdLLzilambda11777  zdLLzilambda11777R33 (gzdLLzilambda11777R33[106:7], gzdLLzilambda11777R33[6:0], callResR133);
  assign gzdLLzilambda11777R34 = {gMainzidev[99:0], 7'h22};
  zdLLzilambda11777  zdLLzilambda11777R34 (gzdLLzilambda11777R34[106:7], gzdLLzilambda11777R34[6:0], callResR134);
  assign gzdLLzilambda11777R35 = {gMainzidev[99:0], 7'h23};
  zdLLzilambda11777  zdLLzilambda11777R35 (gzdLLzilambda11777R35[106:7], gzdLLzilambda11777R35[6:0], callResR135);
  assign gzdLLzilambda11777R36 = {gMainzidev[99:0], 7'h24};
  zdLLzilambda11777  zdLLzilambda11777R36 (gzdLLzilambda11777R36[106:7], gzdLLzilambda11777R36[6:0], callResR136);
  assign gzdLLzilambda11777R37 = {gMainzidev[99:0], 7'h25};
  zdLLzilambda11777  zdLLzilambda11777R37 (gzdLLzilambda11777R37[106:7], gzdLLzilambda11777R37[6:0], callResR137);
  assign gzdLLzilambda11777R38 = {gMainzidev[99:0], 7'h26};
  zdLLzilambda11777  zdLLzilambda11777R38 (gzdLLzilambda11777R38[106:7], gzdLLzilambda11777R38[6:0], callResR138);
  assign gzdLLzilambda11777R39 = {gMainzidev[99:0], 7'h27};
  zdLLzilambda11777  zdLLzilambda11777R39 (gzdLLzilambda11777R39[106:7], gzdLLzilambda11777R39[6:0], callResR139);
  assign gzdLLzilambda11777R40 = {gMainzidev[99:0], 7'h28};
  zdLLzilambda11777  zdLLzilambda11777R40 (gzdLLzilambda11777R40[106:7], gzdLLzilambda11777R40[6:0], callResR140);
  assign gzdLLzilambda11777R41 = {gMainzidev[99:0], 7'h29};
  zdLLzilambda11777  zdLLzilambda11777R41 (gzdLLzilambda11777R41[106:7], gzdLLzilambda11777R41[6:0], callResR141);
  assign gzdLLzilambda11777R42 = {gMainzidev[99:0], 7'h2a};
  zdLLzilambda11777  zdLLzilambda11777R42 (gzdLLzilambda11777R42[106:7], gzdLLzilambda11777R42[6:0], callResR142);
  assign gzdLLzilambda11777R43 = {gMainzidev[99:0], 7'h2b};
  zdLLzilambda11777  zdLLzilambda11777R43 (gzdLLzilambda11777R43[106:7], gzdLLzilambda11777R43[6:0], callResR143);
  assign gzdLLzilambda11777R44 = {gMainzidev[99:0], 7'h2c};
  zdLLzilambda11777  zdLLzilambda11777R44 (gzdLLzilambda11777R44[106:7], gzdLLzilambda11777R44[6:0], callResR144);
  assign gzdLLzilambda11777R45 = {gMainzidev[99:0], 7'h2d};
  zdLLzilambda11777  zdLLzilambda11777R45 (gzdLLzilambda11777R45[106:7], gzdLLzilambda11777R45[6:0], callResR145);
  assign gzdLLzilambda11777R46 = {gMainzidev[99:0], 7'h2e};
  zdLLzilambda11777  zdLLzilambda11777R46 (gzdLLzilambda11777R46[106:7], gzdLLzilambda11777R46[6:0], callResR146);
  assign gzdLLzilambda11777R47 = {gMainzidev[99:0], 7'h2f};
  zdLLzilambda11777  zdLLzilambda11777R47 (gzdLLzilambda11777R47[106:7], gzdLLzilambda11777R47[6:0], callResR147);
  assign gzdLLzilambda11777R48 = {gMainzidev[99:0], 7'h30};
  zdLLzilambda11777  zdLLzilambda11777R48 (gzdLLzilambda11777R48[106:7], gzdLLzilambda11777R48[6:0], callResR148);
  assign gzdLLzilambda11777R49 = {gMainzidev[99:0], 7'h31};
  zdLLzilambda11777  zdLLzilambda11777R49 (gzdLLzilambda11777R49[106:7], gzdLLzilambda11777R49[6:0], callResR149);
  assign gzdLLzilambda11777R50 = {gMainzidev[99:0], 7'h32};
  zdLLzilambda11777  zdLLzilambda11777R50 (gzdLLzilambda11777R50[106:7], gzdLLzilambda11777R50[6:0], callResR150);
  assign gzdLLzilambda11777R51 = {gMainzidev[99:0], 7'h33};
  zdLLzilambda11777  zdLLzilambda11777R51 (gzdLLzilambda11777R51[106:7], gzdLLzilambda11777R51[6:0], callResR151);
  assign gzdLLzilambda11777R52 = {gMainzidev[99:0], 7'h34};
  zdLLzilambda11777  zdLLzilambda11777R52 (gzdLLzilambda11777R52[106:7], gzdLLzilambda11777R52[6:0], callResR152);
  assign gzdLLzilambda11777R53 = {gMainzidev[99:0], 7'h35};
  zdLLzilambda11777  zdLLzilambda11777R53 (gzdLLzilambda11777R53[106:7], gzdLLzilambda11777R53[6:0], callResR153);
  assign gzdLLzilambda11777R54 = {gMainzidev[99:0], 7'h36};
  zdLLzilambda11777  zdLLzilambda11777R54 (gzdLLzilambda11777R54[106:7], gzdLLzilambda11777R54[6:0], callResR154);
  assign gzdLLzilambda11777R55 = {gMainzidev[99:0], 7'h37};
  zdLLzilambda11777  zdLLzilambda11777R55 (gzdLLzilambda11777R55[106:7], gzdLLzilambda11777R55[6:0], callResR155);
  assign gzdLLzilambda11777R56 = {gMainzidev[99:0], 7'h38};
  zdLLzilambda11777  zdLLzilambda11777R56 (gzdLLzilambda11777R56[106:7], gzdLLzilambda11777R56[6:0], callResR156);
  assign gzdLLzilambda11777R57 = {gMainzidev[99:0], 7'h39};
  zdLLzilambda11777  zdLLzilambda11777R57 (gzdLLzilambda11777R57[106:7], gzdLLzilambda11777R57[6:0], callResR157);
  assign gzdLLzilambda11777R58 = {gMainzidev[99:0], 7'h3a};
  zdLLzilambda11777  zdLLzilambda11777R58 (gzdLLzilambda11777R58[106:7], gzdLLzilambda11777R58[6:0], callResR158);
  assign gzdLLzilambda11777R59 = {gMainzidev[99:0], 7'h3b};
  zdLLzilambda11777  zdLLzilambda11777R59 (gzdLLzilambda11777R59[106:7], gzdLLzilambda11777R59[6:0], callResR159);
  assign gzdLLzilambda11777R60 = {gMainzidev[99:0], 7'h3c};
  zdLLzilambda11777  zdLLzilambda11777R60 (gzdLLzilambda11777R60[106:7], gzdLLzilambda11777R60[6:0], callResR160);
  assign gzdLLzilambda11777R61 = {gMainzidev[99:0], 7'h3d};
  zdLLzilambda11777  zdLLzilambda11777R61 (gzdLLzilambda11777R61[106:7], gzdLLzilambda11777R61[6:0], callResR161);
  assign gzdLLzilambda11777R62 = {gMainzidev[99:0], 7'h3e};
  zdLLzilambda11777  zdLLzilambda11777R62 (gzdLLzilambda11777R62[106:7], gzdLLzilambda11777R62[6:0], callResR162);
  assign gzdLLzilambda11777R63 = {gMainzidev[99:0], 7'h3f};
  zdLLzilambda11777  zdLLzilambda11777R63 (gzdLLzilambda11777R63[106:7], gzdLLzilambda11777R63[6:0], callResR163);
  assign gzdLLzilambda11777R64 = {gMainzidev[99:0], 7'h40};
  zdLLzilambda11777  zdLLzilambda11777R64 (gzdLLzilambda11777R64[106:7], gzdLLzilambda11777R64[6:0], callResR164);
  assign gzdLLzilambda11777R65 = {gMainzidev[99:0], 7'h41};
  zdLLzilambda11777  zdLLzilambda11777R65 (gzdLLzilambda11777R65[106:7], gzdLLzilambda11777R65[6:0], callResR165);
  assign gzdLLzilambda11777R66 = {gMainzidev[99:0], 7'h42};
  zdLLzilambda11777  zdLLzilambda11777R66 (gzdLLzilambda11777R66[106:7], gzdLLzilambda11777R66[6:0], callResR166);
  assign gzdLLzilambda11777R67 = {gMainzidev[99:0], 7'h43};
  zdLLzilambda11777  zdLLzilambda11777R67 (gzdLLzilambda11777R67[106:7], gzdLLzilambda11777R67[6:0], callResR167);
  assign gzdLLzilambda11777R68 = {gMainzidev[99:0], 7'h44};
  zdLLzilambda11777  zdLLzilambda11777R68 (gzdLLzilambda11777R68[106:7], gzdLLzilambda11777R68[6:0], callResR168);
  assign gzdLLzilambda11777R69 = {gMainzidev[99:0], 7'h45};
  zdLLzilambda11777  zdLLzilambda11777R69 (gzdLLzilambda11777R69[106:7], gzdLLzilambda11777R69[6:0], callResR169);
  assign gzdLLzilambda11777R70 = {gMainzidev[99:0], 7'h46};
  zdLLzilambda11777  zdLLzilambda11777R70 (gzdLLzilambda11777R70[106:7], gzdLLzilambda11777R70[6:0], callResR170);
  assign gzdLLzilambda11777R71 = {gMainzidev[99:0], 7'h47};
  zdLLzilambda11777  zdLLzilambda11777R71 (gzdLLzilambda11777R71[106:7], gzdLLzilambda11777R71[6:0], callResR171);
  assign gzdLLzilambda11777R72 = {gMainzidev[99:0], 7'h48};
  zdLLzilambda11777  zdLLzilambda11777R72 (gzdLLzilambda11777R72[106:7], gzdLLzilambda11777R72[6:0], callResR172);
  assign gzdLLzilambda11777R73 = {gMainzidev[99:0], 7'h49};
  zdLLzilambda11777  zdLLzilambda11777R73 (gzdLLzilambda11777R73[106:7], gzdLLzilambda11777R73[6:0], callResR173);
  assign gzdLLzilambda11777R74 = {gMainzidev[99:0], 7'h4a};
  zdLLzilambda11777  zdLLzilambda11777R74 (gzdLLzilambda11777R74[106:7], gzdLLzilambda11777R74[6:0], callResR174);
  assign gzdLLzilambda11777R75 = {gMainzidev[99:0], 7'h4b};
  zdLLzilambda11777  zdLLzilambda11777R75 (gzdLLzilambda11777R75[106:7], gzdLLzilambda11777R75[6:0], callResR175);
  assign gzdLLzilambda11777R76 = {gMainzidev[99:0], 7'h4c};
  zdLLzilambda11777  zdLLzilambda11777R76 (gzdLLzilambda11777R76[106:7], gzdLLzilambda11777R76[6:0], callResR176);
  assign gzdLLzilambda11777R77 = {gMainzidev[99:0], 7'h4d};
  zdLLzilambda11777  zdLLzilambda11777R77 (gzdLLzilambda11777R77[106:7], gzdLLzilambda11777R77[6:0], callResR177);
  assign gzdLLzilambda11777R78 = {gMainzidev[99:0], 7'h4e};
  zdLLzilambda11777  zdLLzilambda11777R78 (gzdLLzilambda11777R78[106:7], gzdLLzilambda11777R78[6:0], callResR178);
  assign gzdLLzilambda11777R79 = {gMainzidev[99:0], 7'h4f};
  zdLLzilambda11777  zdLLzilambda11777R79 (gzdLLzilambda11777R79[106:7], gzdLLzilambda11777R79[6:0], callResR179);
  assign gzdLLzilambda11777R80 = {gMainzidev[99:0], 7'h50};
  zdLLzilambda11777  zdLLzilambda11777R80 (gzdLLzilambda11777R80[106:7], gzdLLzilambda11777R80[6:0], callResR180);
  assign gzdLLzilambda11777R81 = {gMainzidev[99:0], 7'h51};
  zdLLzilambda11777  zdLLzilambda11777R81 (gzdLLzilambda11777R81[106:7], gzdLLzilambda11777R81[6:0], callResR181);
  assign gzdLLzilambda11777R82 = {gMainzidev[99:0], 7'h52};
  zdLLzilambda11777  zdLLzilambda11777R82 (gzdLLzilambda11777R82[106:7], gzdLLzilambda11777R82[6:0], callResR182);
  assign gzdLLzilambda11777R83 = {gMainzidev[99:0], 7'h53};
  zdLLzilambda11777  zdLLzilambda11777R83 (gzdLLzilambda11777R83[106:7], gzdLLzilambda11777R83[6:0], callResR183);
  assign gzdLLzilambda11777R84 = {gMainzidev[99:0], 7'h54};
  zdLLzilambda11777  zdLLzilambda11777R84 (gzdLLzilambda11777R84[106:7], gzdLLzilambda11777R84[6:0], callResR184);
  assign gzdLLzilambda11777R85 = {gMainzidev[99:0], 7'h55};
  zdLLzilambda11777  zdLLzilambda11777R85 (gzdLLzilambda11777R85[106:7], gzdLLzilambda11777R85[6:0], callResR185);
  assign gzdLLzilambda11777R86 = {gMainzidev[99:0], 7'h56};
  zdLLzilambda11777  zdLLzilambda11777R86 (gzdLLzilambda11777R86[106:7], gzdLLzilambda11777R86[6:0], callResR186);
  assign gzdLLzilambda11777R87 = {gMainzidev[99:0], 7'h57};
  zdLLzilambda11777  zdLLzilambda11777R87 (gzdLLzilambda11777R87[106:7], gzdLLzilambda11777R87[6:0], callResR187);
  assign gzdLLzilambda11777R88 = {gMainzidev[99:0], 7'h58};
  zdLLzilambda11777  zdLLzilambda11777R88 (gzdLLzilambda11777R88[106:7], gzdLLzilambda11777R88[6:0], callResR188);
  assign gzdLLzilambda11777R89 = {gMainzidev[99:0], 7'h59};
  zdLLzilambda11777  zdLLzilambda11777R89 (gzdLLzilambda11777R89[106:7], gzdLLzilambda11777R89[6:0], callResR189);
  assign gzdLLzilambda11777R90 = {gMainzidev[99:0], 7'h5a};
  zdLLzilambda11777  zdLLzilambda11777R90 (gzdLLzilambda11777R90[106:7], gzdLLzilambda11777R90[6:0], callResR190);
  assign gzdLLzilambda11777R91 = {gMainzidev[99:0], 7'h5b};
  zdLLzilambda11777  zdLLzilambda11777R91 (gzdLLzilambda11777R91[106:7], gzdLLzilambda11777R91[6:0], callResR191);
  assign gzdLLzilambda11777R92 = {gMainzidev[99:0], 7'h5c};
  zdLLzilambda11777  zdLLzilambda11777R92 (gzdLLzilambda11777R92[106:7], gzdLLzilambda11777R92[6:0], callResR192);
  assign gzdLLzilambda11777R93 = {gMainzidev[99:0], 7'h5d};
  zdLLzilambda11777  zdLLzilambda11777R93 (gzdLLzilambda11777R93[106:7], gzdLLzilambda11777R93[6:0], callResR193);
  assign gzdLLzilambda11777R94 = {gMainzidev[99:0], 7'h5e};
  zdLLzilambda11777  zdLLzilambda11777R94 (gzdLLzilambda11777R94[106:7], gzdLLzilambda11777R94[6:0], callResR194);
  assign gzdLLzilambda11777R95 = {gMainzidev[99:0], 7'h5f};
  zdLLzilambda11777  zdLLzilambda11777R95 (gzdLLzilambda11777R95[106:7], gzdLLzilambda11777R95[6:0], callResR195);
  assign gzdLLzilambda11777R96 = {gMainzidev[99:0], 7'h60};
  zdLLzilambda11777  zdLLzilambda11777R96 (gzdLLzilambda11777R96[106:7], gzdLLzilambda11777R96[6:0], callResR196);
  assign gzdLLzilambda11777R97 = {gMainzidev[99:0], 7'h61};
  zdLLzilambda11777  zdLLzilambda11777R97 (gzdLLzilambda11777R97[106:7], gzdLLzilambda11777R97[6:0], callResR197);
  assign gzdLLzilambda11777R98 = {gMainzidev[99:0], 7'h62};
  zdLLzilambda11777  zdLLzilambda11777R98 (gzdLLzilambda11777R98[106:7], gzdLLzilambda11777R98[6:0], callResR198);
  assign gzdLLzilambda11777R99 = {gMainzidev[99:0], 7'h63};
  zdLLzilambda11777  zdLLzilambda11777R99 (gzdLLzilambda11777R99[106:7], gzdLLzilambda11777R99[6:0], callResR199);
  assign gzdLLzilambda11786 = {gMainzidev[99:0], 7'h00};
  zdLLzilambda11786  zdLLzilambda11786 (gzdLLzilambda11786[106:7], gzdLLzilambda11786[6:0], callResR200);
  assign gzdLLzilambda11786R1 = {gMainzidev[99:0], 7'h01};
  zdLLzilambda11786  zdLLzilambda11786R1 (gzdLLzilambda11786R1[106:7], gzdLLzilambda11786R1[6:0], callResR201);
  assign gzdLLzilambda11786R2 = {gMainzidev[99:0], 7'h02};
  zdLLzilambda11786  zdLLzilambda11786R2 (gzdLLzilambda11786R2[106:7], gzdLLzilambda11786R2[6:0], callResR202);
  assign gzdLLzilambda11786R3 = {gMainzidev[99:0], 7'h03};
  zdLLzilambda11786  zdLLzilambda11786R3 (gzdLLzilambda11786R3[106:7], gzdLLzilambda11786R3[6:0], callResR203);
  assign gzdLLzilambda11786R4 = {gMainzidev[99:0], 7'h04};
  zdLLzilambda11786  zdLLzilambda11786R4 (gzdLLzilambda11786R4[106:7], gzdLLzilambda11786R4[6:0], callResR204);
  assign gzdLLzilambda11786R5 = {gMainzidev[99:0], 7'h05};
  zdLLzilambda11786  zdLLzilambda11786R5 (gzdLLzilambda11786R5[106:7], gzdLLzilambda11786R5[6:0], callResR205);
  assign gzdLLzilambda11786R6 = {gMainzidev[99:0], 7'h06};
  zdLLzilambda11786  zdLLzilambda11786R6 (gzdLLzilambda11786R6[106:7], gzdLLzilambda11786R6[6:0], callResR206);
  assign gzdLLzilambda11786R7 = {gMainzidev[99:0], 7'h07};
  zdLLzilambda11786  zdLLzilambda11786R7 (gzdLLzilambda11786R7[106:7], gzdLLzilambda11786R7[6:0], callResR207);
  assign gzdLLzilambda11786R8 = {gMainzidev[99:0], 7'h08};
  zdLLzilambda11786  zdLLzilambda11786R8 (gzdLLzilambda11786R8[106:7], gzdLLzilambda11786R8[6:0], callResR208);
  assign gzdLLzilambda11786R9 = {gMainzidev[99:0], 7'h09};
  zdLLzilambda11786  zdLLzilambda11786R9 (gzdLLzilambda11786R9[106:7], gzdLLzilambda11786R9[6:0], callResR209);
  assign gzdLLzilambda11786R10 = {gMainzidev[99:0], 7'h0a};
  zdLLzilambda11786  zdLLzilambda11786R10 (gzdLLzilambda11786R10[106:7], gzdLLzilambda11786R10[6:0], callResR210);
  assign gzdLLzilambda11786R11 = {gMainzidev[99:0], 7'h0b};
  zdLLzilambda11786  zdLLzilambda11786R11 (gzdLLzilambda11786R11[106:7], gzdLLzilambda11786R11[6:0], callResR211);
  assign gzdLLzilambda11786R12 = {gMainzidev[99:0], 7'h0c};
  zdLLzilambda11786  zdLLzilambda11786R12 (gzdLLzilambda11786R12[106:7], gzdLLzilambda11786R12[6:0], callResR212);
  assign gzdLLzilambda11786R13 = {gMainzidev[99:0], 7'h0d};
  zdLLzilambda11786  zdLLzilambda11786R13 (gzdLLzilambda11786R13[106:7], gzdLLzilambda11786R13[6:0], callResR213);
  assign gzdLLzilambda11786R14 = {gMainzidev[99:0], 7'h0e};
  zdLLzilambda11786  zdLLzilambda11786R14 (gzdLLzilambda11786R14[106:7], gzdLLzilambda11786R14[6:0], callResR214);
  assign gzdLLzilambda11786R15 = {gMainzidev[99:0], 7'h0f};
  zdLLzilambda11786  zdLLzilambda11786R15 (gzdLLzilambda11786R15[106:7], gzdLLzilambda11786R15[6:0], callResR215);
  assign gzdLLzilambda11786R16 = {gMainzidev[99:0], 7'h10};
  zdLLzilambda11786  zdLLzilambda11786R16 (gzdLLzilambda11786R16[106:7], gzdLLzilambda11786R16[6:0], callResR216);
  assign gzdLLzilambda11786R17 = {gMainzidev[99:0], 7'h11};
  zdLLzilambda11786  zdLLzilambda11786R17 (gzdLLzilambda11786R17[106:7], gzdLLzilambda11786R17[6:0], callResR217);
  assign gzdLLzilambda11786R18 = {gMainzidev[99:0], 7'h12};
  zdLLzilambda11786  zdLLzilambda11786R18 (gzdLLzilambda11786R18[106:7], gzdLLzilambda11786R18[6:0], callResR218);
  assign gzdLLzilambda11786R19 = {gMainzidev[99:0], 7'h13};
  zdLLzilambda11786  zdLLzilambda11786R19 (gzdLLzilambda11786R19[106:7], gzdLLzilambda11786R19[6:0], callResR219);
  assign gzdLLzilambda11786R20 = {gMainzidev[99:0], 7'h14};
  zdLLzilambda11786  zdLLzilambda11786R20 (gzdLLzilambda11786R20[106:7], gzdLLzilambda11786R20[6:0], callResR220);
  assign gzdLLzilambda11786R21 = {gMainzidev[99:0], 7'h15};
  zdLLzilambda11786  zdLLzilambda11786R21 (gzdLLzilambda11786R21[106:7], gzdLLzilambda11786R21[6:0], callResR221);
  assign gzdLLzilambda11786R22 = {gMainzidev[99:0], 7'h16};
  zdLLzilambda11786  zdLLzilambda11786R22 (gzdLLzilambda11786R22[106:7], gzdLLzilambda11786R22[6:0], callResR222);
  assign gzdLLzilambda11786R23 = {gMainzidev[99:0], 7'h17};
  zdLLzilambda11786  zdLLzilambda11786R23 (gzdLLzilambda11786R23[106:7], gzdLLzilambda11786R23[6:0], callResR223);
  assign gzdLLzilambda11786R24 = {gMainzidev[99:0], 7'h18};
  zdLLzilambda11786  zdLLzilambda11786R24 (gzdLLzilambda11786R24[106:7], gzdLLzilambda11786R24[6:0], callResR224);
  assign gzdLLzilambda11786R25 = {gMainzidev[99:0], 7'h19};
  zdLLzilambda11786  zdLLzilambda11786R25 (gzdLLzilambda11786R25[106:7], gzdLLzilambda11786R25[6:0], callResR225);
  assign gzdLLzilambda11786R26 = {gMainzidev[99:0], 7'h1a};
  zdLLzilambda11786  zdLLzilambda11786R26 (gzdLLzilambda11786R26[106:7], gzdLLzilambda11786R26[6:0], callResR226);
  assign gzdLLzilambda11786R27 = {gMainzidev[99:0], 7'h1b};
  zdLLzilambda11786  zdLLzilambda11786R27 (gzdLLzilambda11786R27[106:7], gzdLLzilambda11786R27[6:0], callResR227);
  assign gzdLLzilambda11786R28 = {gMainzidev[99:0], 7'h1c};
  zdLLzilambda11786  zdLLzilambda11786R28 (gzdLLzilambda11786R28[106:7], gzdLLzilambda11786R28[6:0], callResR228);
  assign gzdLLzilambda11786R29 = {gMainzidev[99:0], 7'h1d};
  zdLLzilambda11786  zdLLzilambda11786R29 (gzdLLzilambda11786R29[106:7], gzdLLzilambda11786R29[6:0], callResR229);
  assign gzdLLzilambda11786R30 = {gMainzidev[99:0], 7'h1e};
  zdLLzilambda11786  zdLLzilambda11786R30 (gzdLLzilambda11786R30[106:7], gzdLLzilambda11786R30[6:0], callResR230);
  assign gzdLLzilambda11786R31 = {gMainzidev[99:0], 7'h1f};
  zdLLzilambda11786  zdLLzilambda11786R31 (gzdLLzilambda11786R31[106:7], gzdLLzilambda11786R31[6:0], callResR231);
  assign gzdLLzilambda11786R32 = {gMainzidev[99:0], 7'h20};
  zdLLzilambda11786  zdLLzilambda11786R32 (gzdLLzilambda11786R32[106:7], gzdLLzilambda11786R32[6:0], callResR232);
  assign gzdLLzilambda11786R33 = {gMainzidev[99:0], 7'h21};
  zdLLzilambda11786  zdLLzilambda11786R33 (gzdLLzilambda11786R33[106:7], gzdLLzilambda11786R33[6:0], callResR233);
  assign gzdLLzilambda11786R34 = {gMainzidev[99:0], 7'h22};
  zdLLzilambda11786  zdLLzilambda11786R34 (gzdLLzilambda11786R34[106:7], gzdLLzilambda11786R34[6:0], callResR234);
  assign gzdLLzilambda11786R35 = {gMainzidev[99:0], 7'h23};
  zdLLzilambda11786  zdLLzilambda11786R35 (gzdLLzilambda11786R35[106:7], gzdLLzilambda11786R35[6:0], callResR235);
  assign gzdLLzilambda11786R36 = {gMainzidev[99:0], 7'h24};
  zdLLzilambda11786  zdLLzilambda11786R36 (gzdLLzilambda11786R36[106:7], gzdLLzilambda11786R36[6:0], callResR236);
  assign gzdLLzilambda11786R37 = {gMainzidev[99:0], 7'h25};
  zdLLzilambda11786  zdLLzilambda11786R37 (gzdLLzilambda11786R37[106:7], gzdLLzilambda11786R37[6:0], callResR237);
  assign gzdLLzilambda11786R38 = {gMainzidev[99:0], 7'h26};
  zdLLzilambda11786  zdLLzilambda11786R38 (gzdLLzilambda11786R38[106:7], gzdLLzilambda11786R38[6:0], callResR238);
  assign gzdLLzilambda11786R39 = {gMainzidev[99:0], 7'h27};
  zdLLzilambda11786  zdLLzilambda11786R39 (gzdLLzilambda11786R39[106:7], gzdLLzilambda11786R39[6:0], callResR239);
  assign gzdLLzilambda11786R40 = {gMainzidev[99:0], 7'h28};
  zdLLzilambda11786  zdLLzilambda11786R40 (gzdLLzilambda11786R40[106:7], gzdLLzilambda11786R40[6:0], callResR240);
  assign gzdLLzilambda11786R41 = {gMainzidev[99:0], 7'h29};
  zdLLzilambda11786  zdLLzilambda11786R41 (gzdLLzilambda11786R41[106:7], gzdLLzilambda11786R41[6:0], callResR241);
  assign gzdLLzilambda11786R42 = {gMainzidev[99:0], 7'h2a};
  zdLLzilambda11786  zdLLzilambda11786R42 (gzdLLzilambda11786R42[106:7], gzdLLzilambda11786R42[6:0], callResR242);
  assign gzdLLzilambda11786R43 = {gMainzidev[99:0], 7'h2b};
  zdLLzilambda11786  zdLLzilambda11786R43 (gzdLLzilambda11786R43[106:7], gzdLLzilambda11786R43[6:0], callResR243);
  assign gzdLLzilambda11786R44 = {gMainzidev[99:0], 7'h2c};
  zdLLzilambda11786  zdLLzilambda11786R44 (gzdLLzilambda11786R44[106:7], gzdLLzilambda11786R44[6:0], callResR244);
  assign gzdLLzilambda11786R45 = {gMainzidev[99:0], 7'h2d};
  zdLLzilambda11786  zdLLzilambda11786R45 (gzdLLzilambda11786R45[106:7], gzdLLzilambda11786R45[6:0], callResR245);
  assign gzdLLzilambda11786R46 = {gMainzidev[99:0], 7'h2e};
  zdLLzilambda11786  zdLLzilambda11786R46 (gzdLLzilambda11786R46[106:7], gzdLLzilambda11786R46[6:0], callResR246);
  assign gzdLLzilambda11786R47 = {gMainzidev[99:0], 7'h2f};
  zdLLzilambda11786  zdLLzilambda11786R47 (gzdLLzilambda11786R47[106:7], gzdLLzilambda11786R47[6:0], callResR247);
  assign gzdLLzilambda11786R48 = {gMainzidev[99:0], 7'h30};
  zdLLzilambda11786  zdLLzilambda11786R48 (gzdLLzilambda11786R48[106:7], gzdLLzilambda11786R48[6:0], callResR248);
  assign gzdLLzilambda11786R49 = {gMainzidev[99:0], 7'h31};
  zdLLzilambda11786  zdLLzilambda11786R49 (gzdLLzilambda11786R49[106:7], gzdLLzilambda11786R49[6:0], callResR249);
  assign gzdLLzilambda11786R50 = {gMainzidev[99:0], 7'h32};
  zdLLzilambda11786  zdLLzilambda11786R50 (gzdLLzilambda11786R50[106:7], gzdLLzilambda11786R50[6:0], callResR250);
  assign gzdLLzilambda11786R51 = {gMainzidev[99:0], 7'h33};
  zdLLzilambda11786  zdLLzilambda11786R51 (gzdLLzilambda11786R51[106:7], gzdLLzilambda11786R51[6:0], callResR251);
  assign gzdLLzilambda11786R52 = {gMainzidev[99:0], 7'h34};
  zdLLzilambda11786  zdLLzilambda11786R52 (gzdLLzilambda11786R52[106:7], gzdLLzilambda11786R52[6:0], callResR252);
  assign gzdLLzilambda11786R53 = {gMainzidev[99:0], 7'h35};
  zdLLzilambda11786  zdLLzilambda11786R53 (gzdLLzilambda11786R53[106:7], gzdLLzilambda11786R53[6:0], callResR253);
  assign gzdLLzilambda11786R54 = {gMainzidev[99:0], 7'h36};
  zdLLzilambda11786  zdLLzilambda11786R54 (gzdLLzilambda11786R54[106:7], gzdLLzilambda11786R54[6:0], callResR254);
  assign gzdLLzilambda11786R55 = {gMainzidev[99:0], 7'h37};
  zdLLzilambda11786  zdLLzilambda11786R55 (gzdLLzilambda11786R55[106:7], gzdLLzilambda11786R55[6:0], callResR255);
  assign gzdLLzilambda11786R56 = {gMainzidev[99:0], 7'h38};
  zdLLzilambda11786  zdLLzilambda11786R56 (gzdLLzilambda11786R56[106:7], gzdLLzilambda11786R56[6:0], callResR256);
  assign gzdLLzilambda11786R57 = {gMainzidev[99:0], 7'h39};
  zdLLzilambda11786  zdLLzilambda11786R57 (gzdLLzilambda11786R57[106:7], gzdLLzilambda11786R57[6:0], callResR257);
  assign gzdLLzilambda11786R58 = {gMainzidev[99:0], 7'h3a};
  zdLLzilambda11786  zdLLzilambda11786R58 (gzdLLzilambda11786R58[106:7], gzdLLzilambda11786R58[6:0], callResR258);
  assign gzdLLzilambda11786R59 = {gMainzidev[99:0], 7'h3b};
  zdLLzilambda11786  zdLLzilambda11786R59 (gzdLLzilambda11786R59[106:7], gzdLLzilambda11786R59[6:0], callResR259);
  assign gzdLLzilambda11786R60 = {gMainzidev[99:0], 7'h3c};
  zdLLzilambda11786  zdLLzilambda11786R60 (gzdLLzilambda11786R60[106:7], gzdLLzilambda11786R60[6:0], callResR260);
  assign gzdLLzilambda11786R61 = {gMainzidev[99:0], 7'h3d};
  zdLLzilambda11786  zdLLzilambda11786R61 (gzdLLzilambda11786R61[106:7], gzdLLzilambda11786R61[6:0], callResR261);
  assign gzdLLzilambda11786R62 = {gMainzidev[99:0], 7'h3e};
  zdLLzilambda11786  zdLLzilambda11786R62 (gzdLLzilambda11786R62[106:7], gzdLLzilambda11786R62[6:0], callResR262);
  assign gzdLLzilambda11786R63 = {gMainzidev[99:0], 7'h3f};
  zdLLzilambda11786  zdLLzilambda11786R63 (gzdLLzilambda11786R63[106:7], gzdLLzilambda11786R63[6:0], callResR263);
  assign gzdLLzilambda11786R64 = {gMainzidev[99:0], 7'h40};
  zdLLzilambda11786  zdLLzilambda11786R64 (gzdLLzilambda11786R64[106:7], gzdLLzilambda11786R64[6:0], callResR264);
  assign gzdLLzilambda11786R65 = {gMainzidev[99:0], 7'h41};
  zdLLzilambda11786  zdLLzilambda11786R65 (gzdLLzilambda11786R65[106:7], gzdLLzilambda11786R65[6:0], callResR265);
  assign gzdLLzilambda11786R66 = {gMainzidev[99:0], 7'h42};
  zdLLzilambda11786  zdLLzilambda11786R66 (gzdLLzilambda11786R66[106:7], gzdLLzilambda11786R66[6:0], callResR266);
  assign gzdLLzilambda11786R67 = {gMainzidev[99:0], 7'h43};
  zdLLzilambda11786  zdLLzilambda11786R67 (gzdLLzilambda11786R67[106:7], gzdLLzilambda11786R67[6:0], callResR267);
  assign gzdLLzilambda11786R68 = {gMainzidev[99:0], 7'h44};
  zdLLzilambda11786  zdLLzilambda11786R68 (gzdLLzilambda11786R68[106:7], gzdLLzilambda11786R68[6:0], callResR268);
  assign gzdLLzilambda11786R69 = {gMainzidev[99:0], 7'h45};
  zdLLzilambda11786  zdLLzilambda11786R69 (gzdLLzilambda11786R69[106:7], gzdLLzilambda11786R69[6:0], callResR269);
  assign gzdLLzilambda11786R70 = {gMainzidev[99:0], 7'h46};
  zdLLzilambda11786  zdLLzilambda11786R70 (gzdLLzilambda11786R70[106:7], gzdLLzilambda11786R70[6:0], callResR270);
  assign gzdLLzilambda11786R71 = {gMainzidev[99:0], 7'h47};
  zdLLzilambda11786  zdLLzilambda11786R71 (gzdLLzilambda11786R71[106:7], gzdLLzilambda11786R71[6:0], callResR271);
  assign gzdLLzilambda11786R72 = {gMainzidev[99:0], 7'h48};
  zdLLzilambda11786  zdLLzilambda11786R72 (gzdLLzilambda11786R72[106:7], gzdLLzilambda11786R72[6:0], callResR272);
  assign gzdLLzilambda11786R73 = {gMainzidev[99:0], 7'h49};
  zdLLzilambda11786  zdLLzilambda11786R73 (gzdLLzilambda11786R73[106:7], gzdLLzilambda11786R73[6:0], callResR273);
  assign gzdLLzilambda11786R74 = {gMainzidev[99:0], 7'h4a};
  zdLLzilambda11786  zdLLzilambda11786R74 (gzdLLzilambda11786R74[106:7], gzdLLzilambda11786R74[6:0], callResR274);
  assign gzdLLzilambda11786R75 = {gMainzidev[99:0], 7'h4b};
  zdLLzilambda11786  zdLLzilambda11786R75 (gzdLLzilambda11786R75[106:7], gzdLLzilambda11786R75[6:0], callResR275);
  assign gzdLLzilambda11786R76 = {gMainzidev[99:0], 7'h4c};
  zdLLzilambda11786  zdLLzilambda11786R76 (gzdLLzilambda11786R76[106:7], gzdLLzilambda11786R76[6:0], callResR276);
  assign gzdLLzilambda11786R77 = {gMainzidev[99:0], 7'h4d};
  zdLLzilambda11786  zdLLzilambda11786R77 (gzdLLzilambda11786R77[106:7], gzdLLzilambda11786R77[6:0], callResR277);
  assign gzdLLzilambda11786R78 = {gMainzidev[99:0], 7'h4e};
  zdLLzilambda11786  zdLLzilambda11786R78 (gzdLLzilambda11786R78[106:7], gzdLLzilambda11786R78[6:0], callResR278);
  assign gzdLLzilambda11786R79 = {gMainzidev[99:0], 7'h4f};
  zdLLzilambda11786  zdLLzilambda11786R79 (gzdLLzilambda11786R79[106:7], gzdLLzilambda11786R79[6:0], callResR279);
  assign gzdLLzilambda11786R80 = {gMainzidev[99:0], 7'h50};
  zdLLzilambda11786  zdLLzilambda11786R80 (gzdLLzilambda11786R80[106:7], gzdLLzilambda11786R80[6:0], callResR280);
  assign gzdLLzilambda11786R81 = {gMainzidev[99:0], 7'h51};
  zdLLzilambda11786  zdLLzilambda11786R81 (gzdLLzilambda11786R81[106:7], gzdLLzilambda11786R81[6:0], callResR281);
  assign gzdLLzilambda11786R82 = {gMainzidev[99:0], 7'h52};
  zdLLzilambda11786  zdLLzilambda11786R82 (gzdLLzilambda11786R82[106:7], gzdLLzilambda11786R82[6:0], callResR282);
  assign gzdLLzilambda11786R83 = {gMainzidev[99:0], 7'h53};
  zdLLzilambda11786  zdLLzilambda11786R83 (gzdLLzilambda11786R83[106:7], gzdLLzilambda11786R83[6:0], callResR283);
  assign gzdLLzilambda11786R84 = {gMainzidev[99:0], 7'h54};
  zdLLzilambda11786  zdLLzilambda11786R84 (gzdLLzilambda11786R84[106:7], gzdLLzilambda11786R84[6:0], callResR284);
  assign gzdLLzilambda11786R85 = {gMainzidev[99:0], 7'h55};
  zdLLzilambda11786  zdLLzilambda11786R85 (gzdLLzilambda11786R85[106:7], gzdLLzilambda11786R85[6:0], callResR285);
  assign gzdLLzilambda11786R86 = {gMainzidev[99:0], 7'h56};
  zdLLzilambda11786  zdLLzilambda11786R86 (gzdLLzilambda11786R86[106:7], gzdLLzilambda11786R86[6:0], callResR286);
  assign gzdLLzilambda11786R87 = {gMainzidev[99:0], 7'h57};
  zdLLzilambda11786  zdLLzilambda11786R87 (gzdLLzilambda11786R87[106:7], gzdLLzilambda11786R87[6:0], callResR287);
  assign gzdLLzilambda11786R88 = {gMainzidev[99:0], 7'h58};
  zdLLzilambda11786  zdLLzilambda11786R88 (gzdLLzilambda11786R88[106:7], gzdLLzilambda11786R88[6:0], callResR288);
  assign gzdLLzilambda11786R89 = {gMainzidev[99:0], 7'h59};
  zdLLzilambda11786  zdLLzilambda11786R89 (gzdLLzilambda11786R89[106:7], gzdLLzilambda11786R89[6:0], callResR289);
  assign gzdLLzilambda11786R90 = {gMainzidev[99:0], 7'h5a};
  zdLLzilambda11786  zdLLzilambda11786R90 (gzdLLzilambda11786R90[106:7], gzdLLzilambda11786R90[6:0], callResR290);
  assign gzdLLzilambda11786R91 = {gMainzidev[99:0], 7'h5b};
  zdLLzilambda11786  zdLLzilambda11786R91 (gzdLLzilambda11786R91[106:7], gzdLLzilambda11786R91[6:0], callResR291);
  assign gzdLLzilambda11786R92 = {gMainzidev[99:0], 7'h5c};
  zdLLzilambda11786  zdLLzilambda11786R92 (gzdLLzilambda11786R92[106:7], gzdLLzilambda11786R92[6:0], callResR292);
  assign gzdLLzilambda11786R93 = {gMainzidev[99:0], 7'h5d};
  zdLLzilambda11786  zdLLzilambda11786R93 (gzdLLzilambda11786R93[106:7], gzdLLzilambda11786R93[6:0], callResR293);
  assign gzdLLzilambda11786R94 = {gMainzidev[99:0], 7'h5e};
  zdLLzilambda11786  zdLLzilambda11786R94 (gzdLLzilambda11786R94[106:7], gzdLLzilambda11786R94[6:0], callResR294);
  assign gzdLLzilambda11786R95 = {gMainzidev[99:0], 7'h5f};
  zdLLzilambda11786  zdLLzilambda11786R95 (gzdLLzilambda11786R95[106:7], gzdLLzilambda11786R95[6:0], callResR295);
  assign gzdLLzilambda11786R96 = {gMainzidev[99:0], 7'h60};
  zdLLzilambda11786  zdLLzilambda11786R96 (gzdLLzilambda11786R96[106:7], gzdLLzilambda11786R96[6:0], callResR296);
  assign gzdLLzilambda11786R97 = {gMainzidev[99:0], 7'h61};
  zdLLzilambda11786  zdLLzilambda11786R97 (gzdLLzilambda11786R97[106:7], gzdLLzilambda11786R97[6:0], callResR297);
  assign gzdLLzilambda11786R98 = {gMainzidev[99:0], 7'h62};
  zdLLzilambda11786  zdLLzilambda11786R98 (gzdLLzilambda11786R98[106:7], gzdLLzilambda11786R98[6:0], callResR298);
  assign gzdLLzilambda11786R99 = {gMainzidev[99:0], 7'h63};
  zdLLzilambda11786  zdLLzilambda11786R99 (gzdLLzilambda11786R99[106:7], gzdLLzilambda11786R99[6:0], callResR299);
  assign gzdLLzilambda11795 = {gMainzidev[99:0], 7'h00};
  zdLLzilambda11795  zdLLzilambda11795 (gzdLLzilambda11795[106:7], gzdLLzilambda11795[6:0], callResR300);
  assign gzdLLzilambda11795R1 = {gMainzidev[99:0], 7'h01};
  zdLLzilambda11795  zdLLzilambda11795R1 (gzdLLzilambda11795R1[106:7], gzdLLzilambda11795R1[6:0], callResR301);
  assign gzdLLzilambda11795R2 = {gMainzidev[99:0], 7'h02};
  zdLLzilambda11795  zdLLzilambda11795R2 (gzdLLzilambda11795R2[106:7], gzdLLzilambda11795R2[6:0], callResR302);
  assign gzdLLzilambda11795R3 = {gMainzidev[99:0], 7'h03};
  zdLLzilambda11795  zdLLzilambda11795R3 (gzdLLzilambda11795R3[106:7], gzdLLzilambda11795R3[6:0], callResR303);
  assign gzdLLzilambda11795R4 = {gMainzidev[99:0], 7'h04};
  zdLLzilambda11795  zdLLzilambda11795R4 (gzdLLzilambda11795R4[106:7], gzdLLzilambda11795R4[6:0], callResR304);
  assign gzdLLzilambda11795R5 = {gMainzidev[99:0], 7'h05};
  zdLLzilambda11795  zdLLzilambda11795R5 (gzdLLzilambda11795R5[106:7], gzdLLzilambda11795R5[6:0], callResR305);
  assign gzdLLzilambda11795R6 = {gMainzidev[99:0], 7'h06};
  zdLLzilambda11795  zdLLzilambda11795R6 (gzdLLzilambda11795R6[106:7], gzdLLzilambda11795R6[6:0], callResR306);
  assign gzdLLzilambda11795R7 = {gMainzidev[99:0], 7'h07};
  zdLLzilambda11795  zdLLzilambda11795R7 (gzdLLzilambda11795R7[106:7], gzdLLzilambda11795R7[6:0], callResR307);
  assign gzdLLzilambda11795R8 = {gMainzidev[99:0], 7'h08};
  zdLLzilambda11795  zdLLzilambda11795R8 (gzdLLzilambda11795R8[106:7], gzdLLzilambda11795R8[6:0], callResR308);
  assign gzdLLzilambda11795R9 = {gMainzidev[99:0], 7'h09};
  zdLLzilambda11795  zdLLzilambda11795R9 (gzdLLzilambda11795R9[106:7], gzdLLzilambda11795R9[6:0], callResR309);
  assign gzdLLzilambda11795R10 = {gMainzidev[99:0], 7'h0a};
  zdLLzilambda11795  zdLLzilambda11795R10 (gzdLLzilambda11795R10[106:7], gzdLLzilambda11795R10[6:0], callResR310);
  assign gzdLLzilambda11795R11 = {gMainzidev[99:0], 7'h0b};
  zdLLzilambda11795  zdLLzilambda11795R11 (gzdLLzilambda11795R11[106:7], gzdLLzilambda11795R11[6:0], callResR311);
  assign gzdLLzilambda11795R12 = {gMainzidev[99:0], 7'h0c};
  zdLLzilambda11795  zdLLzilambda11795R12 (gzdLLzilambda11795R12[106:7], gzdLLzilambda11795R12[6:0], callResR312);
  assign gzdLLzilambda11795R13 = {gMainzidev[99:0], 7'h0d};
  zdLLzilambda11795  zdLLzilambda11795R13 (gzdLLzilambda11795R13[106:7], gzdLLzilambda11795R13[6:0], callResR313);
  assign gzdLLzilambda11795R14 = {gMainzidev[99:0], 7'h0e};
  zdLLzilambda11795  zdLLzilambda11795R14 (gzdLLzilambda11795R14[106:7], gzdLLzilambda11795R14[6:0], callResR314);
  assign gzdLLzilambda11795R15 = {gMainzidev[99:0], 7'h0f};
  zdLLzilambda11795  zdLLzilambda11795R15 (gzdLLzilambda11795R15[106:7], gzdLLzilambda11795R15[6:0], callResR315);
  assign gzdLLzilambda11795R16 = {gMainzidev[99:0], 7'h10};
  zdLLzilambda11795  zdLLzilambda11795R16 (gzdLLzilambda11795R16[106:7], gzdLLzilambda11795R16[6:0], callResR316);
  assign gzdLLzilambda11795R17 = {gMainzidev[99:0], 7'h11};
  zdLLzilambda11795  zdLLzilambda11795R17 (gzdLLzilambda11795R17[106:7], gzdLLzilambda11795R17[6:0], callResR317);
  assign gzdLLzilambda11795R18 = {gMainzidev[99:0], 7'h12};
  zdLLzilambda11795  zdLLzilambda11795R18 (gzdLLzilambda11795R18[106:7], gzdLLzilambda11795R18[6:0], callResR318);
  assign gzdLLzilambda11795R19 = {gMainzidev[99:0], 7'h13};
  zdLLzilambda11795  zdLLzilambda11795R19 (gzdLLzilambda11795R19[106:7], gzdLLzilambda11795R19[6:0], callResR319);
  assign gzdLLzilambda11795R20 = {gMainzidev[99:0], 7'h14};
  zdLLzilambda11795  zdLLzilambda11795R20 (gzdLLzilambda11795R20[106:7], gzdLLzilambda11795R20[6:0], callResR320);
  assign gzdLLzilambda11795R21 = {gMainzidev[99:0], 7'h15};
  zdLLzilambda11795  zdLLzilambda11795R21 (gzdLLzilambda11795R21[106:7], gzdLLzilambda11795R21[6:0], callResR321);
  assign gzdLLzilambda11795R22 = {gMainzidev[99:0], 7'h16};
  zdLLzilambda11795  zdLLzilambda11795R22 (gzdLLzilambda11795R22[106:7], gzdLLzilambda11795R22[6:0], callResR322);
  assign gzdLLzilambda11795R23 = {gMainzidev[99:0], 7'h17};
  zdLLzilambda11795  zdLLzilambda11795R23 (gzdLLzilambda11795R23[106:7], gzdLLzilambda11795R23[6:0], callResR323);
  assign gzdLLzilambda11795R24 = {gMainzidev[99:0], 7'h18};
  zdLLzilambda11795  zdLLzilambda11795R24 (gzdLLzilambda11795R24[106:7], gzdLLzilambda11795R24[6:0], callResR324);
  assign gzdLLzilambda11795R25 = {gMainzidev[99:0], 7'h19};
  zdLLzilambda11795  zdLLzilambda11795R25 (gzdLLzilambda11795R25[106:7], gzdLLzilambda11795R25[6:0], callResR325);
  assign gzdLLzilambda11795R26 = {gMainzidev[99:0], 7'h1a};
  zdLLzilambda11795  zdLLzilambda11795R26 (gzdLLzilambda11795R26[106:7], gzdLLzilambda11795R26[6:0], callResR326);
  assign gzdLLzilambda11795R27 = {gMainzidev[99:0], 7'h1b};
  zdLLzilambda11795  zdLLzilambda11795R27 (gzdLLzilambda11795R27[106:7], gzdLLzilambda11795R27[6:0], callResR327);
  assign gzdLLzilambda11795R28 = {gMainzidev[99:0], 7'h1c};
  zdLLzilambda11795  zdLLzilambda11795R28 (gzdLLzilambda11795R28[106:7], gzdLLzilambda11795R28[6:0], callResR328);
  assign gzdLLzilambda11795R29 = {gMainzidev[99:0], 7'h1d};
  zdLLzilambda11795  zdLLzilambda11795R29 (gzdLLzilambda11795R29[106:7], gzdLLzilambda11795R29[6:0], callResR329);
  assign gzdLLzilambda11795R30 = {gMainzidev[99:0], 7'h1e};
  zdLLzilambda11795  zdLLzilambda11795R30 (gzdLLzilambda11795R30[106:7], gzdLLzilambda11795R30[6:0], callResR330);
  assign gzdLLzilambda11795R31 = {gMainzidev[99:0], 7'h1f};
  zdLLzilambda11795  zdLLzilambda11795R31 (gzdLLzilambda11795R31[106:7], gzdLLzilambda11795R31[6:0], callResR331);
  assign gzdLLzilambda11795R32 = {gMainzidev[99:0], 7'h20};
  zdLLzilambda11795  zdLLzilambda11795R32 (gzdLLzilambda11795R32[106:7], gzdLLzilambda11795R32[6:0], callResR332);
  assign gzdLLzilambda11795R33 = {gMainzidev[99:0], 7'h21};
  zdLLzilambda11795  zdLLzilambda11795R33 (gzdLLzilambda11795R33[106:7], gzdLLzilambda11795R33[6:0], callResR333);
  assign gzdLLzilambda11795R34 = {gMainzidev[99:0], 7'h22};
  zdLLzilambda11795  zdLLzilambda11795R34 (gzdLLzilambda11795R34[106:7], gzdLLzilambda11795R34[6:0], callResR334);
  assign gzdLLzilambda11795R35 = {gMainzidev[99:0], 7'h23};
  zdLLzilambda11795  zdLLzilambda11795R35 (gzdLLzilambda11795R35[106:7], gzdLLzilambda11795R35[6:0], callResR335);
  assign gzdLLzilambda11795R36 = {gMainzidev[99:0], 7'h24};
  zdLLzilambda11795  zdLLzilambda11795R36 (gzdLLzilambda11795R36[106:7], gzdLLzilambda11795R36[6:0], callResR336);
  assign gzdLLzilambda11795R37 = {gMainzidev[99:0], 7'h25};
  zdLLzilambda11795  zdLLzilambda11795R37 (gzdLLzilambda11795R37[106:7], gzdLLzilambda11795R37[6:0], callResR337);
  assign gzdLLzilambda11795R38 = {gMainzidev[99:0], 7'h26};
  zdLLzilambda11795  zdLLzilambda11795R38 (gzdLLzilambda11795R38[106:7], gzdLLzilambda11795R38[6:0], callResR338);
  assign gzdLLzilambda11795R39 = {gMainzidev[99:0], 7'h27};
  zdLLzilambda11795  zdLLzilambda11795R39 (gzdLLzilambda11795R39[106:7], gzdLLzilambda11795R39[6:0], callResR339);
  assign gzdLLzilambda11795R40 = {gMainzidev[99:0], 7'h28};
  zdLLzilambda11795  zdLLzilambda11795R40 (gzdLLzilambda11795R40[106:7], gzdLLzilambda11795R40[6:0], callResR340);
  assign gzdLLzilambda11795R41 = {gMainzidev[99:0], 7'h29};
  zdLLzilambda11795  zdLLzilambda11795R41 (gzdLLzilambda11795R41[106:7], gzdLLzilambda11795R41[6:0], callResR341);
  assign gzdLLzilambda11795R42 = {gMainzidev[99:0], 7'h2a};
  zdLLzilambda11795  zdLLzilambda11795R42 (gzdLLzilambda11795R42[106:7], gzdLLzilambda11795R42[6:0], callResR342);
  assign gzdLLzilambda11795R43 = {gMainzidev[99:0], 7'h2b};
  zdLLzilambda11795  zdLLzilambda11795R43 (gzdLLzilambda11795R43[106:7], gzdLLzilambda11795R43[6:0], callResR343);
  assign gzdLLzilambda11795R44 = {gMainzidev[99:0], 7'h2c};
  zdLLzilambda11795  zdLLzilambda11795R44 (gzdLLzilambda11795R44[106:7], gzdLLzilambda11795R44[6:0], callResR344);
  assign gzdLLzilambda11795R45 = {gMainzidev[99:0], 7'h2d};
  zdLLzilambda11795  zdLLzilambda11795R45 (gzdLLzilambda11795R45[106:7], gzdLLzilambda11795R45[6:0], callResR345);
  assign gzdLLzilambda11795R46 = {gMainzidev[99:0], 7'h2e};
  zdLLzilambda11795  zdLLzilambda11795R46 (gzdLLzilambda11795R46[106:7], gzdLLzilambda11795R46[6:0], callResR346);
  assign gzdLLzilambda11795R47 = {gMainzidev[99:0], 7'h2f};
  zdLLzilambda11795  zdLLzilambda11795R47 (gzdLLzilambda11795R47[106:7], gzdLLzilambda11795R47[6:0], callResR347);
  assign gzdLLzilambda11795R48 = {gMainzidev[99:0], 7'h30};
  zdLLzilambda11795  zdLLzilambda11795R48 (gzdLLzilambda11795R48[106:7], gzdLLzilambda11795R48[6:0], callResR348);
  assign gzdLLzilambda11795R49 = {gMainzidev[99:0], 7'h31};
  zdLLzilambda11795  zdLLzilambda11795R49 (gzdLLzilambda11795R49[106:7], gzdLLzilambda11795R49[6:0], callResR349);
  assign gzdLLzilambda11795R50 = {gMainzidev[99:0], 7'h32};
  zdLLzilambda11795  zdLLzilambda11795R50 (gzdLLzilambda11795R50[106:7], gzdLLzilambda11795R50[6:0], callResR350);
  assign gzdLLzilambda11795R51 = {gMainzidev[99:0], 7'h33};
  zdLLzilambda11795  zdLLzilambda11795R51 (gzdLLzilambda11795R51[106:7], gzdLLzilambda11795R51[6:0], callResR351);
  assign gzdLLzilambda11795R52 = {gMainzidev[99:0], 7'h34};
  zdLLzilambda11795  zdLLzilambda11795R52 (gzdLLzilambda11795R52[106:7], gzdLLzilambda11795R52[6:0], callResR352);
  assign gzdLLzilambda11795R53 = {gMainzidev[99:0], 7'h35};
  zdLLzilambda11795  zdLLzilambda11795R53 (gzdLLzilambda11795R53[106:7], gzdLLzilambda11795R53[6:0], callResR353);
  assign gzdLLzilambda11795R54 = {gMainzidev[99:0], 7'h36};
  zdLLzilambda11795  zdLLzilambda11795R54 (gzdLLzilambda11795R54[106:7], gzdLLzilambda11795R54[6:0], callResR354);
  assign gzdLLzilambda11795R55 = {gMainzidev[99:0], 7'h37};
  zdLLzilambda11795  zdLLzilambda11795R55 (gzdLLzilambda11795R55[106:7], gzdLLzilambda11795R55[6:0], callResR355);
  assign gzdLLzilambda11795R56 = {gMainzidev[99:0], 7'h38};
  zdLLzilambda11795  zdLLzilambda11795R56 (gzdLLzilambda11795R56[106:7], gzdLLzilambda11795R56[6:0], callResR356);
  assign gzdLLzilambda11795R57 = {gMainzidev[99:0], 7'h39};
  zdLLzilambda11795  zdLLzilambda11795R57 (gzdLLzilambda11795R57[106:7], gzdLLzilambda11795R57[6:0], callResR357);
  assign gzdLLzilambda11795R58 = {gMainzidev[99:0], 7'h3a};
  zdLLzilambda11795  zdLLzilambda11795R58 (gzdLLzilambda11795R58[106:7], gzdLLzilambda11795R58[6:0], callResR358);
  assign gzdLLzilambda11795R59 = {gMainzidev[99:0], 7'h3b};
  zdLLzilambda11795  zdLLzilambda11795R59 (gzdLLzilambda11795R59[106:7], gzdLLzilambda11795R59[6:0], callResR359);
  assign gzdLLzilambda11795R60 = {gMainzidev[99:0], 7'h3c};
  zdLLzilambda11795  zdLLzilambda11795R60 (gzdLLzilambda11795R60[106:7], gzdLLzilambda11795R60[6:0], callResR360);
  assign gzdLLzilambda11795R61 = {gMainzidev[99:0], 7'h3d};
  zdLLzilambda11795  zdLLzilambda11795R61 (gzdLLzilambda11795R61[106:7], gzdLLzilambda11795R61[6:0], callResR361);
  assign gzdLLzilambda11795R62 = {gMainzidev[99:0], 7'h3e};
  zdLLzilambda11795  zdLLzilambda11795R62 (gzdLLzilambda11795R62[106:7], gzdLLzilambda11795R62[6:0], callResR362);
  assign gzdLLzilambda11795R63 = {gMainzidev[99:0], 7'h3f};
  zdLLzilambda11795  zdLLzilambda11795R63 (gzdLLzilambda11795R63[106:7], gzdLLzilambda11795R63[6:0], callResR363);
  assign gzdLLzilambda11795R64 = {gMainzidev[99:0], 7'h40};
  zdLLzilambda11795  zdLLzilambda11795R64 (gzdLLzilambda11795R64[106:7], gzdLLzilambda11795R64[6:0], callResR364);
  assign gzdLLzilambda11795R65 = {gMainzidev[99:0], 7'h41};
  zdLLzilambda11795  zdLLzilambda11795R65 (gzdLLzilambda11795R65[106:7], gzdLLzilambda11795R65[6:0], callResR365);
  assign gzdLLzilambda11795R66 = {gMainzidev[99:0], 7'h42};
  zdLLzilambda11795  zdLLzilambda11795R66 (gzdLLzilambda11795R66[106:7], gzdLLzilambda11795R66[6:0], callResR366);
  assign gzdLLzilambda11795R67 = {gMainzidev[99:0], 7'h43};
  zdLLzilambda11795  zdLLzilambda11795R67 (gzdLLzilambda11795R67[106:7], gzdLLzilambda11795R67[6:0], callResR367);
  assign gzdLLzilambda11795R68 = {gMainzidev[99:0], 7'h44};
  zdLLzilambda11795  zdLLzilambda11795R68 (gzdLLzilambda11795R68[106:7], gzdLLzilambda11795R68[6:0], callResR368);
  assign gzdLLzilambda11795R69 = {gMainzidev[99:0], 7'h45};
  zdLLzilambda11795  zdLLzilambda11795R69 (gzdLLzilambda11795R69[106:7], gzdLLzilambda11795R69[6:0], callResR369);
  assign gzdLLzilambda11795R70 = {gMainzidev[99:0], 7'h46};
  zdLLzilambda11795  zdLLzilambda11795R70 (gzdLLzilambda11795R70[106:7], gzdLLzilambda11795R70[6:0], callResR370);
  assign gzdLLzilambda11795R71 = {gMainzidev[99:0], 7'h47};
  zdLLzilambda11795  zdLLzilambda11795R71 (gzdLLzilambda11795R71[106:7], gzdLLzilambda11795R71[6:0], callResR371);
  assign gzdLLzilambda11795R72 = {gMainzidev[99:0], 7'h48};
  zdLLzilambda11795  zdLLzilambda11795R72 (gzdLLzilambda11795R72[106:7], gzdLLzilambda11795R72[6:0], callResR372);
  assign gzdLLzilambda11795R73 = {gMainzidev[99:0], 7'h49};
  zdLLzilambda11795  zdLLzilambda11795R73 (gzdLLzilambda11795R73[106:7], gzdLLzilambda11795R73[6:0], callResR373);
  assign gzdLLzilambda11795R74 = {gMainzidev[99:0], 7'h4a};
  zdLLzilambda11795  zdLLzilambda11795R74 (gzdLLzilambda11795R74[106:7], gzdLLzilambda11795R74[6:0], callResR374);
  assign gzdLLzilambda11795R75 = {gMainzidev[99:0], 7'h4b};
  zdLLzilambda11795  zdLLzilambda11795R75 (gzdLLzilambda11795R75[106:7], gzdLLzilambda11795R75[6:0], callResR375);
  assign gzdLLzilambda11795R76 = {gMainzidev[99:0], 7'h4c};
  zdLLzilambda11795  zdLLzilambda11795R76 (gzdLLzilambda11795R76[106:7], gzdLLzilambda11795R76[6:0], callResR376);
  assign gzdLLzilambda11795R77 = {gMainzidev[99:0], 7'h4d};
  zdLLzilambda11795  zdLLzilambda11795R77 (gzdLLzilambda11795R77[106:7], gzdLLzilambda11795R77[6:0], callResR377);
  assign gzdLLzilambda11795R78 = {gMainzidev[99:0], 7'h4e};
  zdLLzilambda11795  zdLLzilambda11795R78 (gzdLLzilambda11795R78[106:7], gzdLLzilambda11795R78[6:0], callResR378);
  assign gzdLLzilambda11795R79 = {gMainzidev[99:0], 7'h4f};
  zdLLzilambda11795  zdLLzilambda11795R79 (gzdLLzilambda11795R79[106:7], gzdLLzilambda11795R79[6:0], callResR379);
  assign gzdLLzilambda11795R80 = {gMainzidev[99:0], 7'h50};
  zdLLzilambda11795  zdLLzilambda11795R80 (gzdLLzilambda11795R80[106:7], gzdLLzilambda11795R80[6:0], callResR380);
  assign gzdLLzilambda11795R81 = {gMainzidev[99:0], 7'h51};
  zdLLzilambda11795  zdLLzilambda11795R81 (gzdLLzilambda11795R81[106:7], gzdLLzilambda11795R81[6:0], callResR381);
  assign gzdLLzilambda11795R82 = {gMainzidev[99:0], 7'h52};
  zdLLzilambda11795  zdLLzilambda11795R82 (gzdLLzilambda11795R82[106:7], gzdLLzilambda11795R82[6:0], callResR382);
  assign gzdLLzilambda11795R83 = {gMainzidev[99:0], 7'h53};
  zdLLzilambda11795  zdLLzilambda11795R83 (gzdLLzilambda11795R83[106:7], gzdLLzilambda11795R83[6:0], callResR383);
  assign gzdLLzilambda11795R84 = {gMainzidev[99:0], 7'h54};
  zdLLzilambda11795  zdLLzilambda11795R84 (gzdLLzilambda11795R84[106:7], gzdLLzilambda11795R84[6:0], callResR384);
  assign gzdLLzilambda11795R85 = {gMainzidev[99:0], 7'h55};
  zdLLzilambda11795  zdLLzilambda11795R85 (gzdLLzilambda11795R85[106:7], gzdLLzilambda11795R85[6:0], callResR385);
  assign gzdLLzilambda11795R86 = {gMainzidev[99:0], 7'h56};
  zdLLzilambda11795  zdLLzilambda11795R86 (gzdLLzilambda11795R86[106:7], gzdLLzilambda11795R86[6:0], callResR386);
  assign gzdLLzilambda11795R87 = {gMainzidev[99:0], 7'h57};
  zdLLzilambda11795  zdLLzilambda11795R87 (gzdLLzilambda11795R87[106:7], gzdLLzilambda11795R87[6:0], callResR387);
  assign gzdLLzilambda11795R88 = {gMainzidev[99:0], 7'h58};
  zdLLzilambda11795  zdLLzilambda11795R88 (gzdLLzilambda11795R88[106:7], gzdLLzilambda11795R88[6:0], callResR388);
  assign gzdLLzilambda11795R89 = {gMainzidev[99:0], 7'h59};
  zdLLzilambda11795  zdLLzilambda11795R89 (gzdLLzilambda11795R89[106:7], gzdLLzilambda11795R89[6:0], callResR389);
  assign gzdLLzilambda11795R90 = {gMainzidev[99:0], 7'h5a};
  zdLLzilambda11795  zdLLzilambda11795R90 (gzdLLzilambda11795R90[106:7], gzdLLzilambda11795R90[6:0], callResR390);
  assign gzdLLzilambda11795R91 = {gMainzidev[99:0], 7'h5b};
  zdLLzilambda11795  zdLLzilambda11795R91 (gzdLLzilambda11795R91[106:7], gzdLLzilambda11795R91[6:0], callResR391);
  assign gzdLLzilambda11795R92 = {gMainzidev[99:0], 7'h5c};
  zdLLzilambda11795  zdLLzilambda11795R92 (gzdLLzilambda11795R92[106:7], gzdLLzilambda11795R92[6:0], callResR392);
  assign gzdLLzilambda11795R93 = {gMainzidev[99:0], 7'h5d};
  zdLLzilambda11795  zdLLzilambda11795R93 (gzdLLzilambda11795R93[106:7], gzdLLzilambda11795R93[6:0], callResR393);
  assign gzdLLzilambda11795R94 = {gMainzidev[99:0], 7'h5e};
  zdLLzilambda11795  zdLLzilambda11795R94 (gzdLLzilambda11795R94[106:7], gzdLLzilambda11795R94[6:0], callResR394);
  assign gzdLLzilambda11795R95 = {gMainzidev[99:0], 7'h5f};
  zdLLzilambda11795  zdLLzilambda11795R95 (gzdLLzilambda11795R95[106:7], gzdLLzilambda11795R95[6:0], callResR395);
  assign gzdLLzilambda11795R96 = {gMainzidev[99:0], 7'h60};
  zdLLzilambda11795  zdLLzilambda11795R96 (gzdLLzilambda11795R96[106:7], gzdLLzilambda11795R96[6:0], callResR396);
  assign gzdLLzilambda11795R97 = {gMainzidev[99:0], 7'h61};
  zdLLzilambda11795  zdLLzilambda11795R97 (gzdLLzilambda11795R97[106:7], gzdLLzilambda11795R97[6:0], callResR397);
  assign gzdLLzilambda11795R98 = {gMainzidev[99:0], 7'h62};
  zdLLzilambda11795  zdLLzilambda11795R98 (gzdLLzilambda11795R98[106:7], gzdLLzilambda11795R98[6:0], callResR398);
  assign gzdLLzilambda11795R99 = {gMainzidev[99:0], 7'h63};
  zdLLzilambda11795  zdLLzilambda11795R99 (gzdLLzilambda11795R99[106:7], gzdLLzilambda11795R99[6:0], callResR399);
  assign res = {1'h1, callRes, callResR1, callResR2, callResR3, callResR4, callResR5, callResR6, callResR7, callResR8, callResR9, callResR10, callResR11, callResR12, callResR13, callResR14, callResR15, callResR16, callResR17, callResR18, callResR19, callResR20, callResR21, callResR22, callResR23, callResR24, callResR25, callResR26, callResR27, callResR28, callResR29, callResR30, callResR31, callResR32, callResR33, callResR34, callResR35, callResR36, callResR37, callResR38, callResR39, callResR40, callResR41, callResR42, callResR43, callResR44, callResR45, callResR46, callResR47, callResR48, callResR49, callResR50, callResR51, callResR52, callResR53, callResR54, callResR55, callResR56, callResR57, callResR58, callResR59, callResR60, callResR61, callResR62, callResR63, callResR64, callResR65, callResR66, callResR67, callResR68, callResR69, callResR70, callResR71, callResR72, callResR73, callResR74, callResR75, callResR76, callResR77, callResR78, callResR79, callResR80, callResR81, callResR82, callResR83, callResR84, callResR85, callResR86, callResR87, callResR88, callResR89, callResR90, callResR91, callResR92, callResR93, callResR94, callResR95, callResR96, callResR97, callResR98, callResR99, callResR100, callResR101, callResR102, callResR103, callResR104, callResR105, callResR106, callResR107, callResR108, callResR109, callResR110, callResR111, callResR112, callResR113, callResR114, callResR115, callResR116, callResR117, callResR118, callResR119, callResR120, callResR121, callResR122, callResR123, callResR124, callResR125, callResR126, callResR127, callResR128, callResR129, callResR130, callResR131, callResR132, callResR133, callResR134, callResR135, callResR136, callResR137, callResR138, callResR139, callResR140, callResR141, callResR142, callResR143, callResR144, callResR145, callResR146, callResR147, callResR148, callResR149, callResR150, callResR151, callResR152, callResR153, callResR154, callResR155, callResR156, callResR157, callResR158, callResR159, callResR160, callResR161, callResR162, callResR163, callResR164, callResR165, callResR166, callResR167, callResR168, callResR169, callResR170, callResR171, callResR172, callResR173, callResR174, callResR175, callResR176, callResR177, callResR178, callResR179, callResR180, callResR181, callResR182, callResR183, callResR184, callResR185, callResR186, callResR187, callResR188, callResR189, callResR190, callResR191, callResR192, callResR193, callResR194, callResR195, callResR196, callResR197, callResR198, callResR199, callResR200, callResR201, callResR202, callResR203, callResR204, callResR205, callResR206, callResR207, callResR208, callResR209, callResR210, callResR211, callResR212, callResR213, callResR214, callResR215, callResR216, callResR217, callResR218, callResR219, callResR220, callResR221, callResR222, callResR223, callResR224, callResR225, callResR226, callResR227, callResR228, callResR229, callResR230, callResR231, callResR232, callResR233, callResR234, callResR235, callResR236, callResR237, callResR238, callResR239, callResR240, callResR241, callResR242, callResR243, callResR244, callResR245, callResR246, callResR247, callResR248, callResR249, callResR250, callResR251, callResR252, callResR253, callResR254, callResR255, callResR256, callResR257, callResR258, callResR259, callResR260, callResR261, callResR262, callResR263, callResR264, callResR265, callResR266, callResR267, callResR268, callResR269, callResR270, callResR271, callResR272, callResR273, callResR274, callResR275, callResR276, callResR277, callResR278, callResR279, callResR280, callResR281, callResR282, callResR283, callResR284, callResR285, callResR286, callResR287, callResR288, callResR289, callResR290, callResR291, callResR292, callResR293, callResR294, callResR295, callResR296, callResR297, callResR298, callResR299, callResR300, callResR301, callResR302, callResR303, callResR304, callResR305, callResR306, callResR307, callResR308, callResR309, callResR310, callResR311, callResR312, callResR313, callResR314, callResR315, callResR316, callResR317, callResR318, callResR319, callResR320, callResR321, callResR322, callResR323, callResR324, callResR325, callResR326, callResR327, callResR328, callResR329, callResR330, callResR331, callResR332, callResR333, callResR334, callResR335, callResR336, callResR337, callResR338, callResR339, callResR340, callResR341, callResR342, callResR343, callResR344, callResR345, callResR346, callResR347, callResR348, callResR349, callResR350, callResR351, callResR352, callResR353, callResR354, callResR355, callResR356, callResR357, callResR358, callResR359, callResR360, callResR361, callResR362, callResR363, callResR364, callResR365, callResR366, callResR367, callResR368, callResR369, callResR370, callResR371, callResR372, callResR373, callResR374, callResR375, callResR376, callResR377, callResR378, callResR379, callResR380, callResR381, callResR382, callResR383, callResR384, callResR385, callResR386, callResR387, callResR388, callResR389, callResR390, callResR391, callResR392, callResR393, callResR394, callResR395, callResR396, callResR397, callResR398, callResR399, 1'h0};
endmodule

module zdLLzilambda11768 (input logic [99:0] arg0,
  input logic [6:0] arg1,
  output logic [0:0] res);
  logic [6:0] resizze;
  logic [127:0] resizzeR1;
  logic [0:0] msbit;
  logic [0:0] gReWireziPreludezinot;
  logic [0:0] callRes;
  logic [6:0] resizzeR2;
  logic [127:0] resizzeR3;
  logic [0:0] msbitR1;
  logic [0:0] gReWireziPreludezinotR1;
  logic [0:0] callResR1;
  logic [107:0] gzdLLzicase11762;
  logic [99:0] gMainzix2;
  logic [99:0] callResR2;
  logic [99:0] resizzeR4;
  logic [6:0] resizzeR5;
  logic [255:0] binOp;
  logic [255:0] binOpR1;
  logic [127:0] resizzeR6;
  logic [6:0] resizzeR7;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR8;
  logic [6:0] resizzeR9;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [127:0] resizzeR10;
  logic [107:0] gzdLLzicase11765;
  logic [99:0] resizzeR11;
  logic [6:0] resizzeR12;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [127:0] resizzeR13;
  logic [6:0] resizzeR14;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [127:0] resizzeR15;
  assign resizze = arg1;
  assign resizzeR1 = 128'(resizze[6:0]);
  assign msbit = resizzeR1[0];
  assign gReWireziPreludezinot = msbit[0];
  ReWireziPreludezinot  ReWireziPreludezinot (gReWireziPreludezinot[0], callRes);
  assign resizzeR2 = arg1;
  assign resizzeR3 = 128'(resizzeR2[6:0]);
  assign msbitR1 = resizzeR3[0];
  assign gReWireziPreludezinotR1 = msbitR1[0];
  ReWireziPreludezinot  ReWireziPreludezinotR1 (gReWireziPreludezinotR1[0], callResR1);
  assign gzdLLzicase11762 = {callResR1, arg0, arg1};
  assign gMainzix2 = gzdLLzicase11762[106:7];
  Mainzix2  Mainzix2 (gMainzix2[99:0], callResR2);
  assign resizzeR4 = callResR2;
  assign resizzeR5 = gzdLLzicase11762[6:0];
  assign binOp = {128'(resizzeR5[6:0]), 128'h00000000000000000000000000000001};
  assign binOpR1 = {binOp[255:128] - binOp[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR6 = binOpR1[255:128] % binOpR1[127:0];
  assign resizzeR7 = resizzeR6[6:0];
  assign binOpR2 = {128'(resizzeR7[6:0]), 128'h00000000000000000000000000000002};
  assign binOpR3 = {binOpR2[255:128] / binOpR2[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR8 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR9 = resizzeR8[6:0];
  assign binOpR4 = {128'h00000000000000000000000000000064, 128'(resizzeR9[6:0])};
  assign binOpR5 = {binOpR4[255:128] - binOpR4[127:0], 128'h00000000000000000000000000000001};
  assign binOpR6 = {binOpR5[255:128] - binOpR5[127:0], 128'h00000000000000000000000000000001};
  assign binOpR7 = {128'(resizzeR4[99:0]), binOpR6[255:128] * binOpR6[127:0]};
  assign resizzeR10 = binOpR7[255:128] >> binOpR7[127:0];
  assign gzdLLzicase11765 = {callRes, arg0, arg1};
  assign resizzeR11 = gzdLLzicase11765[106:7];
  assign resizzeR12 = gzdLLzicase11765[6:0];
  assign binOpR8 = {128'(resizzeR12[6:0]), 128'h00000000000000000000000000000002};
  assign binOpR9 = {binOpR8[255:128] / binOpR8[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR13 = binOpR9[255:128] % binOpR9[127:0];
  assign resizzeR14 = resizzeR13[6:0];
  assign binOpR10 = {128'h00000000000000000000000000000064, 128'(resizzeR14[6:0])};
  assign binOpR11 = {binOpR10[255:128] - binOpR10[127:0], 128'h00000000000000000000000000000001};
  assign binOpR12 = {binOpR11[255:128] - binOpR11[127:0], 128'h00000000000000000000000000000001};
  assign binOpR13 = {128'(resizzeR11[99:0]), binOpR12[255:128] * binOpR12[127:0]};
  assign resizzeR15 = binOpR13[255:128] >> binOpR13[127:0];
  assign res = (gzdLLzicase11765[107] == 1'h1) ? resizzeR15[0] : resizzeR10[0];
endmodule

module zdLLzilambda11777 (input logic [99:0] arg0,
  input logic [6:0] arg1,
  output logic [0:0] res);
  logic [6:0] resizze;
  logic [127:0] resizzeR1;
  logic [0:0] msbit;
  logic [0:0] gReWireziPreludezinot;
  logic [0:0] callRes;
  logic [6:0] resizzeR2;
  logic [127:0] resizzeR3;
  logic [0:0] msbitR1;
  logic [0:0] gReWireziPreludezinotR1;
  logic [0:0] callResR1;
  logic [107:0] gzdLLzicase11771;
  logic [99:0] gMainzix2;
  logic [99:0] callResR2;
  logic [99:0] resizzeR4;
  logic [6:0] resizzeR5;
  logic [255:0] binOp;
  logic [255:0] binOpR1;
  logic [127:0] resizzeR6;
  logic [6:0] resizzeR7;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR8;
  logic [6:0] resizzeR9;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR10;
  logic [6:0] resizzeR11;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [127:0] resizzeR12;
  logic [107:0] gzdLLzicase11774;
  logic [99:0] resizzeR13;
  logic [6:0] resizzeR14;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [127:0] resizzeR15;
  logic [6:0] resizzeR16;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [127:0] resizzeR17;
  logic [6:0] resizzeR18;
  logic [255:0] binOpR14;
  logic [255:0] binOpR15;
  logic [255:0] binOpR16;
  logic [255:0] binOpR17;
  logic [127:0] resizzeR19;
  assign resizze = arg1;
  assign resizzeR1 = 128'(resizze[6:0]);
  assign msbit = resizzeR1[0];
  assign gReWireziPreludezinot = msbit[0];
  ReWireziPreludezinot  ReWireziPreludezinot (gReWireziPreludezinot[0], callRes);
  assign resizzeR2 = arg1;
  assign resizzeR3 = 128'(resizzeR2[6:0]);
  assign msbitR1 = resizzeR3[0];
  assign gReWireziPreludezinotR1 = msbitR1[0];
  ReWireziPreludezinot  ReWireziPreludezinotR1 (gReWireziPreludezinotR1[0], callResR1);
  assign gzdLLzicase11771 = {callResR1, arg0, arg1};
  assign gMainzix2 = gzdLLzicase11771[106:7];
  Mainzix2  Mainzix2 (gMainzix2[99:0], callResR2);
  assign resizzeR4 = callResR2;
  assign resizzeR5 = gzdLLzicase11771[6:0];
  assign binOp = {128'(resizzeR5[6:0]), 128'h00000000000000000000000000000001};
  assign binOpR1 = {binOp[255:128] - binOp[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR6 = binOpR1[255:128] % binOpR1[127:0];
  assign resizzeR7 = resizzeR6[6:0];
  assign binOpR2 = {128'h00000000000000000000000000000031, 128'(resizzeR7[6:0])};
  assign binOpR3 = {binOpR2[255:128] + binOpR2[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR8 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR9 = resizzeR8[6:0];
  assign binOpR4 = {128'(resizzeR9[6:0]), 128'h00000000000000000000000000000002};
  assign binOpR5 = {binOpR4[255:128] / binOpR4[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR10 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR11 = resizzeR10[6:0];
  assign binOpR6 = {128'h00000000000000000000000000000064, 128'(resizzeR11[6:0])};
  assign binOpR7 = {binOpR6[255:128] - binOpR6[127:0], 128'h00000000000000000000000000000001};
  assign binOpR8 = {binOpR7[255:128] - binOpR7[127:0], 128'h00000000000000000000000000000001};
  assign binOpR9 = {128'(resizzeR4[99:0]), binOpR8[255:128] * binOpR8[127:0]};
  assign resizzeR12 = binOpR9[255:128] >> binOpR9[127:0];
  assign gzdLLzicase11774 = {callRes, arg0, arg1};
  assign resizzeR13 = gzdLLzicase11774[106:7];
  assign resizzeR14 = gzdLLzicase11774[6:0];
  assign binOpR10 = {128'h00000000000000000000000000000031, 128'(resizzeR14[6:0])};
  assign binOpR11 = {binOpR10[255:128] + binOpR10[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR15 = binOpR11[255:128] % binOpR11[127:0];
  assign resizzeR16 = resizzeR15[6:0];
  assign binOpR12 = {128'(resizzeR16[6:0]), 128'h00000000000000000000000000000002};
  assign binOpR13 = {binOpR12[255:128] / binOpR12[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR17 = binOpR13[255:128] % binOpR13[127:0];
  assign resizzeR18 = resizzeR17[6:0];
  assign binOpR14 = {128'h00000000000000000000000000000064, 128'(resizzeR18[6:0])};
  assign binOpR15 = {binOpR14[255:128] - binOpR14[127:0], 128'h00000000000000000000000000000001};
  assign binOpR16 = {binOpR15[255:128] - binOpR15[127:0], 128'h00000000000000000000000000000001};
  assign binOpR17 = {128'(resizzeR13[99:0]), binOpR16[255:128] * binOpR16[127:0]};
  assign resizzeR19 = binOpR17[255:128] >> binOpR17[127:0];
  assign res = (gzdLLzicase11774[107] == 1'h1) ? resizzeR19[0] : resizzeR12[0];
endmodule

module zdLLzilambda11786 (input logic [99:0] arg0,
  input logic [6:0] arg1,
  output logic [0:0] res);
  logic [6:0] resizze;
  logic [255:0] binOp;
  logic [6:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [107:0] gzdLLzicase11780;
  logic [99:0] gMainzix2;
  logic [99:0] callRes;
  logic [99:0] resizzeR2;
  logic [6:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [6:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR6;
  logic [6:0] resizzeR7;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [127:0] resizzeR8;
  logic [107:0] gzdLLzicase11783;
  logic [99:0] resizzeR9;
  logic [6:0] resizzeR10;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [127:0] resizzeR11;
  logic [6:0] resizzeR12;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [255:0] binOpR14;
  logic [255:0] binOpR15;
  logic [127:0] resizzeR13;
  assign resizze = arg1;
  assign binOp = {128'(resizze[6:0]), 128'h00000000000000000000000000000031};
  assign resizzeR1 = arg1;
  assign binOpR1 = {128'(resizzeR1[6:0]), 128'h00000000000000000000000000000031};
  assign gzdLLzicase11780 = {binOpR1[255:128] < binOpR1[127:0], arg0, arg1};
  assign gMainzix2 = gzdLLzicase11780[106:7];
  Mainzix2  Mainzix2 (gMainzix2[99:0], callRes);
  assign resizzeR2 = callRes;
  assign resizzeR3 = gzdLLzicase11780[6:0];
  assign binOpR2 = {128'(resizzeR3[6:0]), 128'h00000000000000000000000000000031};
  assign binOpR3 = {binOpR2[255:128] - binOpR2[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[6:0];
  assign binOpR4 = {128'(resizzeR5[6:0]), 128'h00000000000000000000000000000002};
  assign binOpR5 = {binOpR4[255:128] * binOpR4[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR6 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR7 = resizzeR6[6:0];
  assign binOpR6 = {128'h00000000000000000000000000000064, 128'(resizzeR7[6:0])};
  assign binOpR7 = {binOpR6[255:128] - binOpR6[127:0], 128'h00000000000000000000000000000001};
  assign binOpR8 = {binOpR7[255:128] - binOpR7[127:0], 128'h00000000000000000000000000000001};
  assign binOpR9 = {128'(resizzeR2[99:0]), binOpR8[255:128] * binOpR8[127:0]};
  assign resizzeR8 = binOpR9[255:128] >> binOpR9[127:0];
  assign gzdLLzicase11783 = {binOp[255:128] < binOp[127:0], arg0, arg1};
  assign resizzeR9 = gzdLLzicase11783[106:7];
  assign resizzeR10 = gzdLLzicase11783[6:0];
  assign binOpR10 = {128'(resizzeR10[6:0]), 128'h00000000000000000000000000000002};
  assign binOpR11 = {binOpR10[255:128] * binOpR10[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR11 = binOpR11[255:128] % binOpR11[127:0];
  assign resizzeR12 = resizzeR11[6:0];
  assign binOpR12 = {128'h00000000000000000000000000000064, 128'(resizzeR12[6:0])};
  assign binOpR13 = {binOpR12[255:128] - binOpR12[127:0], 128'h00000000000000000000000000000001};
  assign binOpR14 = {binOpR13[255:128] - binOpR13[127:0], 128'h00000000000000000000000000000001};
  assign binOpR15 = {128'(resizzeR9[99:0]), binOpR14[255:128] * binOpR14[127:0]};
  assign resizzeR13 = binOpR15[255:128] >> binOpR15[127:0];
  assign res = (gzdLLzicase11783[107] == 1'h1) ? resizzeR13[0] : resizzeR8[0];
endmodule

module zdLLzilambda11795 (input logic [99:0] arg0,
  input logic [6:0] arg1,
  output logic [0:0] res);
  logic [6:0] resizze;
  logic [255:0] binOp;
  logic [6:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [107:0] gzdLLzicase11789;
  logic [99:0] gMainzix2;
  logic [99:0] callRes;
  logic [99:0] resizzeR2;
  logic [6:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [6:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR6;
  logic [6:0] resizzeR7;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [127:0] resizzeR8;
  logic [6:0] resizzeR9;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [127:0] resizzeR10;
  logic [107:0] gzdLLzicase11792;
  logic [99:0] resizzeR11;
  logic [6:0] resizzeR12;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [127:0] resizzeR13;
  logic [6:0] resizzeR14;
  logic [255:0] binOpR14;
  logic [255:0] binOpR15;
  logic [127:0] resizzeR15;
  logic [6:0] resizzeR16;
  logic [255:0] binOpR16;
  logic [255:0] binOpR17;
  logic [255:0] binOpR18;
  logic [255:0] binOpR19;
  logic [127:0] resizzeR17;
  assign resizze = arg1;
  assign binOp = {128'(resizze[6:0]), 128'h00000000000000000000000000000031};
  assign resizzeR1 = arg1;
  assign binOpR1 = {128'(resizzeR1[6:0]), 128'h00000000000000000000000000000031};
  assign gzdLLzicase11789 = {binOpR1[255:128] < binOpR1[127:0], arg0, arg1};
  assign gMainzix2 = gzdLLzicase11789[106:7];
  Mainzix2  Mainzix2 (gMainzix2[99:0], callRes);
  assign resizzeR2 = callRes;
  assign resizzeR3 = gzdLLzicase11789[6:0];
  assign binOpR2 = {128'(resizzeR3[6:0]), 128'h00000000000000000000000000000031};
  assign binOpR3 = {binOpR2[255:128] - binOpR2[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[6:0];
  assign binOpR4 = {128'(resizzeR5[6:0]), 128'h00000000000000000000000000000002};
  assign binOpR5 = {binOpR4[255:128] * binOpR4[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR6 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR7 = resizzeR6[6:0];
  assign binOpR6 = {128'(resizzeR7[6:0]), 128'h00000000000000000000000000000001};
  assign binOpR7 = {binOpR6[255:128] + binOpR6[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR8 = binOpR7[255:128] % binOpR7[127:0];
  assign resizzeR9 = resizzeR8[6:0];
  assign binOpR8 = {128'h00000000000000000000000000000064, 128'(resizzeR9[6:0])};
  assign binOpR9 = {binOpR8[255:128] - binOpR8[127:0], 128'h00000000000000000000000000000001};
  assign binOpR10 = {binOpR9[255:128] - binOpR9[127:0], 128'h00000000000000000000000000000001};
  assign binOpR11 = {128'(resizzeR2[99:0]), binOpR10[255:128] * binOpR10[127:0]};
  assign resizzeR10 = binOpR11[255:128] >> binOpR11[127:0];
  assign gzdLLzicase11792 = {binOp[255:128] < binOp[127:0], arg0, arg1};
  assign resizzeR11 = gzdLLzicase11792[106:7];
  assign resizzeR12 = gzdLLzicase11792[6:0];
  assign binOpR12 = {128'(resizzeR12[6:0]), 128'h00000000000000000000000000000002};
  assign binOpR13 = {binOpR12[255:128] * binOpR12[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR13 = binOpR13[255:128] % binOpR13[127:0];
  assign resizzeR14 = resizzeR13[6:0];
  assign binOpR14 = {128'(resizzeR14[6:0]), 128'h00000000000000000000000000000001};
  assign binOpR15 = {binOpR14[255:128] + binOpR14[127:0], 128'h00000000000000000000000000000064};
  assign resizzeR15 = binOpR15[255:128] % binOpR15[127:0];
  assign resizzeR16 = resizzeR15[6:0];
  assign binOpR16 = {128'h00000000000000000000000000000064, 128'(resizzeR16[6:0])};
  assign binOpR17 = {binOpR16[255:128] - binOpR16[127:0], 128'h00000000000000000000000000000001};
  assign binOpR18 = {binOpR17[255:128] - binOpR17[127:0], 128'h00000000000000000000000000000001};
  assign binOpR19 = {128'(resizzeR11[99:0]), binOpR18[255:128] * binOpR18[127:0]};
  assign resizzeR17 = binOpR19[255:128] >> binOpR19[127:0];
  assign res = (gzdLLzicase11792[107] == 1'h1) ? resizzeR17[0] : resizzeR10[0];
endmodule

module Mainzix2 (input logic [99:0] arg0,
  output logic [99:0] res);
  logic [199:0] binOp;
  assign binOp = {arg0, 100'h0000000000000000000000002};
  assign res = binOp[199:100] * binOp[99:0];
endmodule

module ReWireziPreludezinot (input logic [0:0] arg0,
  output logic [0:0] res);
  logic [0:0] lit;
  assign lit = arg0;
  assign res = (lit[0] == 1'h1) ? 1'h0 : 1'h1;
endmodule