module top_level ();
  logic [0:0] __padding;
  assign __padding = 1'h1;
endmodule