module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [0:0] __in0,
  output logic [1023:0] __out0);
  logic [1024:0] main_nopipeline_in;
  logic [1025:0] zll_main_nopipeline11_in;
  logic [1024:0] zll_main_nopipeline17_in;
  logic [1024:0] zll_main_nopipeline24_in;
  logic [2049:0] zll_main_nopipeline24_out;
  logic [1024:0] zll_main_nopipeline18_in;
  logic [1023:0] zll_main_nopipeline_in;
  logic [2047:0] zll_main_nopipeline15_in;
  logic [2047:0] zll_main_nopipeline19_in;
  logic [1023:0] main_round_in;
  logic [1023:0] zll_main_swap4_in;
  logic [1028:0] main_swapix4_in;
  logic [31:0] main_swapix4_out;
  logic [1028:0] main_swapix4_inR1;
  logic [31:0] main_swapix4_outR1;
  logic [1028:0] main_swapix4_inR2;
  logic [31:0] main_swapix4_outR2;
  logic [1028:0] main_swapix4_inR3;
  logic [31:0] main_swapix4_outR3;
  logic [1028:0] main_swapix4_inR4;
  logic [31:0] main_swapix4_outR4;
  logic [1028:0] main_swapix4_inR5;
  logic [31:0] main_swapix4_outR5;
  logic [1028:0] main_swapix4_inR6;
  logic [31:0] main_swapix4_outR6;
  logic [1028:0] main_swapix4_inR7;
  logic [31:0] main_swapix4_outR7;
  logic [1028:0] main_swapix4_inR8;
  logic [31:0] main_swapix4_outR8;
  logic [1028:0] main_swapix4_inR9;
  logic [31:0] main_swapix4_outR9;
  logic [1028:0] main_swapix4_inR10;
  logic [31:0] main_swapix4_outR10;
  logic [1028:0] main_swapix4_inR11;
  logic [31:0] main_swapix4_outR11;
  logic [1028:0] main_swapix4_inR12;
  logic [31:0] main_swapix4_outR12;
  logic [1028:0] main_swapix4_inR13;
  logic [31:0] main_swapix4_outR13;
  logic [1028:0] main_swapix4_inR14;
  logic [31:0] main_swapix4_outR14;
  logic [1028:0] main_swapix4_inR15;
  logic [31:0] main_swapix4_outR15;
  logic [1028:0] main_swapix4_inR16;
  logic [31:0] main_swapix4_outR16;
  logic [1028:0] main_swapix4_inR17;
  logic [31:0] main_swapix4_outR17;
  logic [1028:0] main_swapix4_inR18;
  logic [31:0] main_swapix4_outR18;
  logic [1028:0] main_swapix4_inR19;
  logic [31:0] main_swapix4_outR19;
  logic [1028:0] main_swapix4_inR20;
  logic [31:0] main_swapix4_outR20;
  logic [1028:0] main_swapix4_inR21;
  logic [31:0] main_swapix4_outR21;
  logic [1028:0] main_swapix4_inR22;
  logic [31:0] main_swapix4_outR22;
  logic [1028:0] main_swapix4_inR23;
  logic [31:0] main_swapix4_outR23;
  logic [1028:0] main_swapix4_inR24;
  logic [31:0] main_swapix4_outR24;
  logic [1028:0] main_swapix4_inR25;
  logic [31:0] main_swapix4_outR25;
  logic [1028:0] main_swapix4_inR26;
  logic [31:0] main_swapix4_outR26;
  logic [1028:0] main_swapix4_inR27;
  logic [31:0] main_swapix4_outR27;
  logic [1028:0] main_swapix4_inR28;
  logic [31:0] main_swapix4_outR28;
  logic [1028:0] main_swapix4_inR29;
  logic [31:0] main_swapix4_outR29;
  logic [1028:0] main_swapix4_inR30;
  logic [31:0] main_swapix4_outR30;
  logic [1028:0] main_swapix4_inR31;
  logic [31:0] main_swapix4_outR31;
  logic [1023:0] zll_main_xor_in;
  logic [1023:0] zll_main_xor_out;
  logic [1023:0] zll_main_swap3_in;
  logic [1028:0] main_swapix3_in;
  logic [31:0] main_swapix3_out;
  logic [1028:0] main_swapix3_inR1;
  logic [31:0] main_swapix3_outR1;
  logic [1028:0] main_swapix3_inR2;
  logic [31:0] main_swapix3_outR2;
  logic [1028:0] main_swapix3_inR3;
  logic [31:0] main_swapix3_outR3;
  logic [1028:0] main_swapix3_inR4;
  logic [31:0] main_swapix3_outR4;
  logic [1028:0] main_swapix3_inR5;
  logic [31:0] main_swapix3_outR5;
  logic [1028:0] main_swapix3_inR6;
  logic [31:0] main_swapix3_outR6;
  logic [1028:0] main_swapix3_inR7;
  logic [31:0] main_swapix3_outR7;
  logic [1028:0] main_swapix3_inR8;
  logic [31:0] main_swapix3_outR8;
  logic [1028:0] main_swapix3_inR9;
  logic [31:0] main_swapix3_outR9;
  logic [1028:0] main_swapix3_inR10;
  logic [31:0] main_swapix3_outR10;
  logic [1028:0] main_swapix3_inR11;
  logic [31:0] main_swapix3_outR11;
  logic [1028:0] main_swapix3_inR12;
  logic [31:0] main_swapix3_outR12;
  logic [1028:0] main_swapix3_inR13;
  logic [31:0] main_swapix3_outR13;
  logic [1028:0] main_swapix3_inR14;
  logic [31:0] main_swapix3_outR14;
  logic [1028:0] main_swapix3_inR15;
  logic [31:0] main_swapix3_outR15;
  logic [1028:0] main_swapix3_inR16;
  logic [31:0] main_swapix3_outR16;
  logic [1028:0] main_swapix3_inR17;
  logic [31:0] main_swapix3_outR17;
  logic [1028:0] main_swapix3_inR18;
  logic [31:0] main_swapix3_outR18;
  logic [1028:0] main_swapix3_inR19;
  logic [31:0] main_swapix3_outR19;
  logic [1028:0] main_swapix3_inR20;
  logic [31:0] main_swapix3_outR20;
  logic [1028:0] main_swapix3_inR21;
  logic [31:0] main_swapix3_outR21;
  logic [1028:0] main_swapix3_inR22;
  logic [31:0] main_swapix3_outR22;
  logic [1028:0] main_swapix3_inR23;
  logic [31:0] main_swapix3_outR23;
  logic [1028:0] main_swapix3_inR24;
  logic [31:0] main_swapix3_outR24;
  logic [1028:0] main_swapix3_inR25;
  logic [31:0] main_swapix3_outR25;
  logic [1028:0] main_swapix3_inR26;
  logic [31:0] main_swapix3_outR26;
  logic [1028:0] main_swapix3_inR27;
  logic [31:0] main_swapix3_outR27;
  logic [1028:0] main_swapix3_inR28;
  logic [31:0] main_swapix3_outR28;
  logic [1028:0] main_swapix3_inR29;
  logic [31:0] main_swapix3_outR29;
  logic [1028:0] main_swapix3_inR30;
  logic [31:0] main_swapix3_outR30;
  logic [1028:0] main_swapix3_inR31;
  logic [31:0] main_swapix3_outR31;
  logic [1023:0] main_rotate_in;
  logic [1055:0] zll_main_rotate_in;
  logic [1023:0] zll_main_rotate_out;
  logic [1023:0] zll_main_add_in;
  logic [1023:0] zll_main_add_out;
  logic [1023:0] zll_main_swap2_in;
  logic [1028:0] main_swapix2_in;
  logic [31:0] main_swapix2_out;
  logic [1028:0] main_swapix2_inR1;
  logic [31:0] main_swapix2_outR1;
  logic [1028:0] main_swapix2_inR2;
  logic [31:0] main_swapix2_outR2;
  logic [1028:0] main_swapix2_inR3;
  logic [31:0] main_swapix2_outR3;
  logic [1028:0] main_swapix2_inR4;
  logic [31:0] main_swapix2_outR4;
  logic [1028:0] main_swapix2_inR5;
  logic [31:0] main_swapix2_outR5;
  logic [1028:0] main_swapix2_inR6;
  logic [31:0] main_swapix2_outR6;
  logic [1028:0] main_swapix2_inR7;
  logic [31:0] main_swapix2_outR7;
  logic [1028:0] main_swapix2_inR8;
  logic [31:0] main_swapix2_outR8;
  logic [1028:0] main_swapix2_inR9;
  logic [31:0] main_swapix2_outR9;
  logic [1028:0] main_swapix2_inR10;
  logic [31:0] main_swapix2_outR10;
  logic [1028:0] main_swapix2_inR11;
  logic [31:0] main_swapix2_outR11;
  logic [1028:0] main_swapix2_inR12;
  logic [31:0] main_swapix2_outR12;
  logic [1028:0] main_swapix2_inR13;
  logic [31:0] main_swapix2_outR13;
  logic [1028:0] main_swapix2_inR14;
  logic [31:0] main_swapix2_outR14;
  logic [1028:0] main_swapix2_inR15;
  logic [31:0] main_swapix2_outR15;
  logic [1028:0] main_swapix2_inR16;
  logic [31:0] main_swapix2_outR16;
  logic [1028:0] main_swapix2_inR17;
  logic [31:0] main_swapix2_outR17;
  logic [1028:0] main_swapix2_inR18;
  logic [31:0] main_swapix2_outR18;
  logic [1028:0] main_swapix2_inR19;
  logic [31:0] main_swapix2_outR19;
  logic [1028:0] main_swapix2_inR20;
  logic [31:0] main_swapix2_outR20;
  logic [1028:0] main_swapix2_inR21;
  logic [31:0] main_swapix2_outR21;
  logic [1028:0] main_swapix2_inR22;
  logic [31:0] main_swapix2_outR22;
  logic [1028:0] main_swapix2_inR23;
  logic [31:0] main_swapix2_outR23;
  logic [1028:0] main_swapix2_inR24;
  logic [31:0] main_swapix2_outR24;
  logic [1028:0] main_swapix2_inR25;
  logic [31:0] main_swapix2_outR25;
  logic [1028:0] main_swapix2_inR26;
  logic [31:0] main_swapix2_outR26;
  logic [1028:0] main_swapix2_inR27;
  logic [31:0] main_swapix2_outR27;
  logic [1028:0] main_swapix2_inR28;
  logic [31:0] main_swapix2_outR28;
  logic [1028:0] main_swapix2_inR29;
  logic [31:0] main_swapix2_outR29;
  logic [1028:0] main_swapix2_inR30;
  logic [31:0] main_swapix2_outR30;
  logic [1028:0] main_swapix2_inR31;
  logic [31:0] main_swapix2_outR31;
  logic [1023:0] zll_main_xor_inR1;
  logic [1023:0] zll_main_xor_outR1;
  logic [1023:0] zll_main_swap1_in;
  logic [1028:0] main_swapix1_in;
  logic [31:0] main_swapix1_out;
  logic [1028:0] main_swapix1_inR1;
  logic [31:0] main_swapix1_outR1;
  logic [1028:0] main_swapix1_inR2;
  logic [31:0] main_swapix1_outR2;
  logic [1028:0] main_swapix1_inR3;
  logic [31:0] main_swapix1_outR3;
  logic [1028:0] main_swapix1_inR4;
  logic [31:0] main_swapix1_outR4;
  logic [1028:0] main_swapix1_inR5;
  logic [31:0] main_swapix1_outR5;
  logic [1028:0] main_swapix1_inR6;
  logic [31:0] main_swapix1_outR6;
  logic [1028:0] main_swapix1_inR7;
  logic [31:0] main_swapix1_outR7;
  logic [1028:0] main_swapix1_inR8;
  logic [31:0] main_swapix1_outR8;
  logic [1028:0] main_swapix1_inR9;
  logic [31:0] main_swapix1_outR9;
  logic [1028:0] main_swapix1_inR10;
  logic [31:0] main_swapix1_outR10;
  logic [1028:0] main_swapix1_inR11;
  logic [31:0] main_swapix1_outR11;
  logic [1028:0] main_swapix1_inR12;
  logic [31:0] main_swapix1_outR12;
  logic [1028:0] main_swapix1_inR13;
  logic [31:0] main_swapix1_outR13;
  logic [1028:0] main_swapix1_inR14;
  logic [31:0] main_swapix1_outR14;
  logic [1028:0] main_swapix1_inR15;
  logic [31:0] main_swapix1_outR15;
  logic [1028:0] main_swapix1_inR16;
  logic [31:0] main_swapix1_outR16;
  logic [1028:0] main_swapix1_inR17;
  logic [31:0] main_swapix1_outR17;
  logic [1028:0] main_swapix1_inR18;
  logic [31:0] main_swapix1_outR18;
  logic [1028:0] main_swapix1_inR19;
  logic [31:0] main_swapix1_outR19;
  logic [1028:0] main_swapix1_inR20;
  logic [31:0] main_swapix1_outR20;
  logic [1028:0] main_swapix1_inR21;
  logic [31:0] main_swapix1_outR21;
  logic [1028:0] main_swapix1_inR22;
  logic [31:0] main_swapix1_outR22;
  logic [1028:0] main_swapix1_inR23;
  logic [31:0] main_swapix1_outR23;
  logic [1028:0] main_swapix1_inR24;
  logic [31:0] main_swapix1_outR24;
  logic [1028:0] main_swapix1_inR25;
  logic [31:0] main_swapix1_outR25;
  logic [1028:0] main_swapix1_inR26;
  logic [31:0] main_swapix1_outR26;
  logic [1028:0] main_swapix1_inR27;
  logic [31:0] main_swapix1_outR27;
  logic [1028:0] main_swapix1_inR28;
  logic [31:0] main_swapix1_outR28;
  logic [1028:0] main_swapix1_inR29;
  logic [31:0] main_swapix1_outR29;
  logic [1028:0] main_swapix1_inR30;
  logic [31:0] main_swapix1_outR30;
  logic [1028:0] main_swapix1_inR31;
  logic [31:0] main_swapix1_outR31;
  logic [1023:0] main_rotate1_in;
  logic [1055:0] zll_main_rotate_inR1;
  logic [1023:0] zll_main_rotate_outR1;
  logic [1023:0] zll_main_add_inR1;
  logic [1023:0] zll_main_add_outR1;
  logic [1023:0] zll_main_nopipeline2_in;
  logic [2049:0] zll_main_nopipeline6_in;
  logic [2049:0] zll_main_nopipeline24_inR1;
  logic [2049:0] zll_main_nopipeline24_outR1;
  logic [1:0] __padding;
  logic [1023:0] __st0;
  logic [1023:0] __st0_next;
  assign main_nopipeline_in = {__in0, __st0};
  assign zll_main_nopipeline11_in = {main_nopipeline_in[1024], main_nopipeline_in[1024], main_nopipeline_in[1023:0]};
  assign zll_main_nopipeline17_in = {zll_main_nopipeline11_in[1025], zll_main_nopipeline11_in[1023:0]};
  assign zll_main_nopipeline24_in = {zll_main_nopipeline17_in[1023:0], zll_main_nopipeline17_in[1024]};
  ZLL_Main_nopipeline24  inst (zll_main_nopipeline24_in[1024:1], zll_main_nopipeline24_out);
  assign zll_main_nopipeline18_in = {zll_main_nopipeline11_in[1023:0], zll_main_nopipeline11_in[1024]};
  assign zll_main_nopipeline_in = zll_main_nopipeline18_in[1024:1];
  assign zll_main_nopipeline15_in = {zll_main_nopipeline_in[1023:0], zll_main_nopipeline_in[1023:0]};
  assign zll_main_nopipeline19_in = zll_main_nopipeline15_in[2047:0];
  assign main_round_in = zll_main_nopipeline19_in[2047:1024];
  assign zll_main_swap4_in = main_round_in[1023:0];
  assign main_swapix4_in = {zll_main_swap4_in[1023:0], 5'h0};
  Main_swapix4  instR1 (main_swapix4_in[1028:5], main_swapix4_in[4:0], main_swapix4_out);
  assign main_swapix4_inR1 = {zll_main_swap4_in[1023:0], 5'h1};
  Main_swapix4  instR2 (main_swapix4_inR1[1028:5], main_swapix4_inR1[4:0], main_swapix4_outR1);
  assign main_swapix4_inR2 = {zll_main_swap4_in[1023:0], 5'h2};
  Main_swapix4  instR3 (main_swapix4_inR2[1028:5], main_swapix4_inR2[4:0], main_swapix4_outR2);
  assign main_swapix4_inR3 = {zll_main_swap4_in[1023:0], 5'h3};
  Main_swapix4  instR4 (main_swapix4_inR3[1028:5], main_swapix4_inR3[4:0], main_swapix4_outR3);
  assign main_swapix4_inR4 = {zll_main_swap4_in[1023:0], 5'h4};
  Main_swapix4  instR5 (main_swapix4_inR4[1028:5], main_swapix4_inR4[4:0], main_swapix4_outR4);
  assign main_swapix4_inR5 = {zll_main_swap4_in[1023:0], 5'h5};
  Main_swapix4  instR6 (main_swapix4_inR5[1028:5], main_swapix4_inR5[4:0], main_swapix4_outR5);
  assign main_swapix4_inR6 = {zll_main_swap4_in[1023:0], 5'h6};
  Main_swapix4  instR7 (main_swapix4_inR6[1028:5], main_swapix4_inR6[4:0], main_swapix4_outR6);
  assign main_swapix4_inR7 = {zll_main_swap4_in[1023:0], 5'h7};
  Main_swapix4  instR8 (main_swapix4_inR7[1028:5], main_swapix4_inR7[4:0], main_swapix4_outR7);
  assign main_swapix4_inR8 = {zll_main_swap4_in[1023:0], 5'h8};
  Main_swapix4  instR9 (main_swapix4_inR8[1028:5], main_swapix4_inR8[4:0], main_swapix4_outR8);
  assign main_swapix4_inR9 = {zll_main_swap4_in[1023:0], 5'h9};
  Main_swapix4  instR10 (main_swapix4_inR9[1028:5], main_swapix4_inR9[4:0], main_swapix4_outR9);
  assign main_swapix4_inR10 = {zll_main_swap4_in[1023:0], 5'ha};
  Main_swapix4  instR11 (main_swapix4_inR10[1028:5], main_swapix4_inR10[4:0], main_swapix4_outR10);
  assign main_swapix4_inR11 = {zll_main_swap4_in[1023:0], 5'hb};
  Main_swapix4  instR12 (main_swapix4_inR11[1028:5], main_swapix4_inR11[4:0], main_swapix4_outR11);
  assign main_swapix4_inR12 = {zll_main_swap4_in[1023:0], 5'hc};
  Main_swapix4  instR13 (main_swapix4_inR12[1028:5], main_swapix4_inR12[4:0], main_swapix4_outR12);
  assign main_swapix4_inR13 = {zll_main_swap4_in[1023:0], 5'hd};
  Main_swapix4  instR14 (main_swapix4_inR13[1028:5], main_swapix4_inR13[4:0], main_swapix4_outR13);
  assign main_swapix4_inR14 = {zll_main_swap4_in[1023:0], 5'he};
  Main_swapix4  instR15 (main_swapix4_inR14[1028:5], main_swapix4_inR14[4:0], main_swapix4_outR14);
  assign main_swapix4_inR15 = {zll_main_swap4_in[1023:0], 5'hf};
  Main_swapix4  instR16 (main_swapix4_inR15[1028:5], main_swapix4_inR15[4:0], main_swapix4_outR15);
  assign main_swapix4_inR16 = {zll_main_swap4_in[1023:0], 5'h10};
  Main_swapix4  instR17 (main_swapix4_inR16[1028:5], main_swapix4_inR16[4:0], main_swapix4_outR16);
  assign main_swapix4_inR17 = {zll_main_swap4_in[1023:0], 5'h11};
  Main_swapix4  instR18 (main_swapix4_inR17[1028:5], main_swapix4_inR17[4:0], main_swapix4_outR17);
  assign main_swapix4_inR18 = {zll_main_swap4_in[1023:0], 5'h12};
  Main_swapix4  instR19 (main_swapix4_inR18[1028:5], main_swapix4_inR18[4:0], main_swapix4_outR18);
  assign main_swapix4_inR19 = {zll_main_swap4_in[1023:0], 5'h13};
  Main_swapix4  instR20 (main_swapix4_inR19[1028:5], main_swapix4_inR19[4:0], main_swapix4_outR19);
  assign main_swapix4_inR20 = {zll_main_swap4_in[1023:0], 5'h14};
  Main_swapix4  instR21 (main_swapix4_inR20[1028:5], main_swapix4_inR20[4:0], main_swapix4_outR20);
  assign main_swapix4_inR21 = {zll_main_swap4_in[1023:0], 5'h15};
  Main_swapix4  instR22 (main_swapix4_inR21[1028:5], main_swapix4_inR21[4:0], main_swapix4_outR21);
  assign main_swapix4_inR22 = {zll_main_swap4_in[1023:0], 5'h16};
  Main_swapix4  instR23 (main_swapix4_inR22[1028:5], main_swapix4_inR22[4:0], main_swapix4_outR22);
  assign main_swapix4_inR23 = {zll_main_swap4_in[1023:0], 5'h17};
  Main_swapix4  instR24 (main_swapix4_inR23[1028:5], main_swapix4_inR23[4:0], main_swapix4_outR23);
  assign main_swapix4_inR24 = {zll_main_swap4_in[1023:0], 5'h18};
  Main_swapix4  instR25 (main_swapix4_inR24[1028:5], main_swapix4_inR24[4:0], main_swapix4_outR24);
  assign main_swapix4_inR25 = {zll_main_swap4_in[1023:0], 5'h19};
  Main_swapix4  instR26 (main_swapix4_inR25[1028:5], main_swapix4_inR25[4:0], main_swapix4_outR25);
  assign main_swapix4_inR26 = {zll_main_swap4_in[1023:0], 5'h1a};
  Main_swapix4  instR27 (main_swapix4_inR26[1028:5], main_swapix4_inR26[4:0], main_swapix4_outR26);
  assign main_swapix4_inR27 = {zll_main_swap4_in[1023:0], 5'h1b};
  Main_swapix4  instR28 (main_swapix4_inR27[1028:5], main_swapix4_inR27[4:0], main_swapix4_outR27);
  assign main_swapix4_inR28 = {zll_main_swap4_in[1023:0], 5'h1c};
  Main_swapix4  instR29 (main_swapix4_inR28[1028:5], main_swapix4_inR28[4:0], main_swapix4_outR28);
  assign main_swapix4_inR29 = {zll_main_swap4_in[1023:0], 5'h1d};
  Main_swapix4  instR30 (main_swapix4_inR29[1028:5], main_swapix4_inR29[4:0], main_swapix4_outR29);
  assign main_swapix4_inR30 = {zll_main_swap4_in[1023:0], 5'h1e};
  Main_swapix4  instR31 (main_swapix4_inR30[1028:5], main_swapix4_inR30[4:0], main_swapix4_outR30);
  assign main_swapix4_inR31 = {zll_main_swap4_in[1023:0], 5'h1f};
  Main_swapix4  instR32 (main_swapix4_inR31[1028:5], main_swapix4_inR31[4:0], main_swapix4_outR31);
  assign zll_main_xor_in = {main_swapix4_out, main_swapix4_outR1, main_swapix4_outR2, main_swapix4_outR3, main_swapix4_outR4, main_swapix4_outR5, main_swapix4_outR6, main_swapix4_outR7, main_swapix4_outR8, main_swapix4_outR9, main_swapix4_outR10, main_swapix4_outR11, main_swapix4_outR12, main_swapix4_outR13, main_swapix4_outR14, main_swapix4_outR15, main_swapix4_outR16, main_swapix4_outR17, main_swapix4_outR18, main_swapix4_outR19, main_swapix4_outR20, main_swapix4_outR21, main_swapix4_outR22, main_swapix4_outR23, main_swapix4_outR24, main_swapix4_outR25, main_swapix4_outR26, main_swapix4_outR27, main_swapix4_outR28, main_swapix4_outR29, main_swapix4_outR30, main_swapix4_outR31};
  ZLL_Main_xor  instR33 (zll_main_xor_in[1023:0], zll_main_xor_out);
  assign zll_main_swap3_in = zll_main_xor_out;
  assign main_swapix3_in = {zll_main_swap3_in[1023:0], 5'h0};
  Main_swapix3  instR34 (main_swapix3_in[1028:5], main_swapix3_in[4:0], main_swapix3_out);
  assign main_swapix3_inR1 = {zll_main_swap3_in[1023:0], 5'h1};
  Main_swapix3  instR35 (main_swapix3_inR1[1028:5], main_swapix3_inR1[4:0], main_swapix3_outR1);
  assign main_swapix3_inR2 = {zll_main_swap3_in[1023:0], 5'h2};
  Main_swapix3  instR36 (main_swapix3_inR2[1028:5], main_swapix3_inR2[4:0], main_swapix3_outR2);
  assign main_swapix3_inR3 = {zll_main_swap3_in[1023:0], 5'h3};
  Main_swapix3  instR37 (main_swapix3_inR3[1028:5], main_swapix3_inR3[4:0], main_swapix3_outR3);
  assign main_swapix3_inR4 = {zll_main_swap3_in[1023:0], 5'h4};
  Main_swapix3  instR38 (main_swapix3_inR4[1028:5], main_swapix3_inR4[4:0], main_swapix3_outR4);
  assign main_swapix3_inR5 = {zll_main_swap3_in[1023:0], 5'h5};
  Main_swapix3  instR39 (main_swapix3_inR5[1028:5], main_swapix3_inR5[4:0], main_swapix3_outR5);
  assign main_swapix3_inR6 = {zll_main_swap3_in[1023:0], 5'h6};
  Main_swapix3  instR40 (main_swapix3_inR6[1028:5], main_swapix3_inR6[4:0], main_swapix3_outR6);
  assign main_swapix3_inR7 = {zll_main_swap3_in[1023:0], 5'h7};
  Main_swapix3  instR41 (main_swapix3_inR7[1028:5], main_swapix3_inR7[4:0], main_swapix3_outR7);
  assign main_swapix3_inR8 = {zll_main_swap3_in[1023:0], 5'h8};
  Main_swapix3  instR42 (main_swapix3_inR8[1028:5], main_swapix3_inR8[4:0], main_swapix3_outR8);
  assign main_swapix3_inR9 = {zll_main_swap3_in[1023:0], 5'h9};
  Main_swapix3  instR43 (main_swapix3_inR9[1028:5], main_swapix3_inR9[4:0], main_swapix3_outR9);
  assign main_swapix3_inR10 = {zll_main_swap3_in[1023:0], 5'ha};
  Main_swapix3  instR44 (main_swapix3_inR10[1028:5], main_swapix3_inR10[4:0], main_swapix3_outR10);
  assign main_swapix3_inR11 = {zll_main_swap3_in[1023:0], 5'hb};
  Main_swapix3  instR45 (main_swapix3_inR11[1028:5], main_swapix3_inR11[4:0], main_swapix3_outR11);
  assign main_swapix3_inR12 = {zll_main_swap3_in[1023:0], 5'hc};
  Main_swapix3  instR46 (main_swapix3_inR12[1028:5], main_swapix3_inR12[4:0], main_swapix3_outR12);
  assign main_swapix3_inR13 = {zll_main_swap3_in[1023:0], 5'hd};
  Main_swapix3  instR47 (main_swapix3_inR13[1028:5], main_swapix3_inR13[4:0], main_swapix3_outR13);
  assign main_swapix3_inR14 = {zll_main_swap3_in[1023:0], 5'he};
  Main_swapix3  instR48 (main_swapix3_inR14[1028:5], main_swapix3_inR14[4:0], main_swapix3_outR14);
  assign main_swapix3_inR15 = {zll_main_swap3_in[1023:0], 5'hf};
  Main_swapix3  instR49 (main_swapix3_inR15[1028:5], main_swapix3_inR15[4:0], main_swapix3_outR15);
  assign main_swapix3_inR16 = {zll_main_swap3_in[1023:0], 5'h10};
  Main_swapix3  instR50 (main_swapix3_inR16[1028:5], main_swapix3_inR16[4:0], main_swapix3_outR16);
  assign main_swapix3_inR17 = {zll_main_swap3_in[1023:0], 5'h11};
  Main_swapix3  instR51 (main_swapix3_inR17[1028:5], main_swapix3_inR17[4:0], main_swapix3_outR17);
  assign main_swapix3_inR18 = {zll_main_swap3_in[1023:0], 5'h12};
  Main_swapix3  instR52 (main_swapix3_inR18[1028:5], main_swapix3_inR18[4:0], main_swapix3_outR18);
  assign main_swapix3_inR19 = {zll_main_swap3_in[1023:0], 5'h13};
  Main_swapix3  instR53 (main_swapix3_inR19[1028:5], main_swapix3_inR19[4:0], main_swapix3_outR19);
  assign main_swapix3_inR20 = {zll_main_swap3_in[1023:0], 5'h14};
  Main_swapix3  instR54 (main_swapix3_inR20[1028:5], main_swapix3_inR20[4:0], main_swapix3_outR20);
  assign main_swapix3_inR21 = {zll_main_swap3_in[1023:0], 5'h15};
  Main_swapix3  instR55 (main_swapix3_inR21[1028:5], main_swapix3_inR21[4:0], main_swapix3_outR21);
  assign main_swapix3_inR22 = {zll_main_swap3_in[1023:0], 5'h16};
  Main_swapix3  instR56 (main_swapix3_inR22[1028:5], main_swapix3_inR22[4:0], main_swapix3_outR22);
  assign main_swapix3_inR23 = {zll_main_swap3_in[1023:0], 5'h17};
  Main_swapix3  instR57 (main_swapix3_inR23[1028:5], main_swapix3_inR23[4:0], main_swapix3_outR23);
  assign main_swapix3_inR24 = {zll_main_swap3_in[1023:0], 5'h18};
  Main_swapix3  instR58 (main_swapix3_inR24[1028:5], main_swapix3_inR24[4:0], main_swapix3_outR24);
  assign main_swapix3_inR25 = {zll_main_swap3_in[1023:0], 5'h19};
  Main_swapix3  instR59 (main_swapix3_inR25[1028:5], main_swapix3_inR25[4:0], main_swapix3_outR25);
  assign main_swapix3_inR26 = {zll_main_swap3_in[1023:0], 5'h1a};
  Main_swapix3  instR60 (main_swapix3_inR26[1028:5], main_swapix3_inR26[4:0], main_swapix3_outR26);
  assign main_swapix3_inR27 = {zll_main_swap3_in[1023:0], 5'h1b};
  Main_swapix3  instR61 (main_swapix3_inR27[1028:5], main_swapix3_inR27[4:0], main_swapix3_outR27);
  assign main_swapix3_inR28 = {zll_main_swap3_in[1023:0], 5'h1c};
  Main_swapix3  instR62 (main_swapix3_inR28[1028:5], main_swapix3_inR28[4:0], main_swapix3_outR28);
  assign main_swapix3_inR29 = {zll_main_swap3_in[1023:0], 5'h1d};
  Main_swapix3  instR63 (main_swapix3_inR29[1028:5], main_swapix3_inR29[4:0], main_swapix3_outR29);
  assign main_swapix3_inR30 = {zll_main_swap3_in[1023:0], 5'h1e};
  Main_swapix3  instR64 (main_swapix3_inR30[1028:5], main_swapix3_inR30[4:0], main_swapix3_outR30);
  assign main_swapix3_inR31 = {zll_main_swap3_in[1023:0], 5'h1f};
  Main_swapix3  instR65 (main_swapix3_inR31[1028:5], main_swapix3_inR31[4:0], main_swapix3_outR31);
  assign main_rotate_in = {main_swapix3_out, main_swapix3_outR1, main_swapix3_outR2, main_swapix3_outR3, main_swapix3_outR4, main_swapix3_outR5, main_swapix3_outR6, main_swapix3_outR7, main_swapix3_outR8, main_swapix3_outR9, main_swapix3_outR10, main_swapix3_outR11, main_swapix3_outR12, main_swapix3_outR13, main_swapix3_outR14, main_swapix3_outR15, main_swapix3_outR16, main_swapix3_outR17, main_swapix3_outR18, main_swapix3_outR19, main_swapix3_outR20, main_swapix3_outR21, main_swapix3_outR22, main_swapix3_outR23, main_swapix3_outR24, main_swapix3_outR25, main_swapix3_outR26, main_swapix3_outR27, main_swapix3_outR28, main_swapix3_outR29, main_swapix3_outR30, main_swapix3_outR31};
  assign zll_main_rotate_in = {32'hb, main_rotate_in[1023:0]};
  ZLL_Main_rotate  instR66 (zll_main_rotate_in[1055:0], zll_main_rotate_out);
  assign zll_main_add_in = zll_main_rotate_out;
  ZLL_Main_add  instR67 (zll_main_add_in[1023:0], zll_main_add_out);
  assign zll_main_swap2_in = zll_main_add_out;
  assign main_swapix2_in = {zll_main_swap2_in[1023:0], 5'h0};
  Main_swapix2  instR68 (main_swapix2_in[1028:5], main_swapix2_in[4:0], main_swapix2_out);
  assign main_swapix2_inR1 = {zll_main_swap2_in[1023:0], 5'h1};
  Main_swapix2  instR69 (main_swapix2_inR1[1028:5], main_swapix2_inR1[4:0], main_swapix2_outR1);
  assign main_swapix2_inR2 = {zll_main_swap2_in[1023:0], 5'h2};
  Main_swapix2  instR70 (main_swapix2_inR2[1028:5], main_swapix2_inR2[4:0], main_swapix2_outR2);
  assign main_swapix2_inR3 = {zll_main_swap2_in[1023:0], 5'h3};
  Main_swapix2  instR71 (main_swapix2_inR3[1028:5], main_swapix2_inR3[4:0], main_swapix2_outR3);
  assign main_swapix2_inR4 = {zll_main_swap2_in[1023:0], 5'h4};
  Main_swapix2  instR72 (main_swapix2_inR4[1028:5], main_swapix2_inR4[4:0], main_swapix2_outR4);
  assign main_swapix2_inR5 = {zll_main_swap2_in[1023:0], 5'h5};
  Main_swapix2  instR73 (main_swapix2_inR5[1028:5], main_swapix2_inR5[4:0], main_swapix2_outR5);
  assign main_swapix2_inR6 = {zll_main_swap2_in[1023:0], 5'h6};
  Main_swapix2  instR74 (main_swapix2_inR6[1028:5], main_swapix2_inR6[4:0], main_swapix2_outR6);
  assign main_swapix2_inR7 = {zll_main_swap2_in[1023:0], 5'h7};
  Main_swapix2  instR75 (main_swapix2_inR7[1028:5], main_swapix2_inR7[4:0], main_swapix2_outR7);
  assign main_swapix2_inR8 = {zll_main_swap2_in[1023:0], 5'h8};
  Main_swapix2  instR76 (main_swapix2_inR8[1028:5], main_swapix2_inR8[4:0], main_swapix2_outR8);
  assign main_swapix2_inR9 = {zll_main_swap2_in[1023:0], 5'h9};
  Main_swapix2  instR77 (main_swapix2_inR9[1028:5], main_swapix2_inR9[4:0], main_swapix2_outR9);
  assign main_swapix2_inR10 = {zll_main_swap2_in[1023:0], 5'ha};
  Main_swapix2  instR78 (main_swapix2_inR10[1028:5], main_swapix2_inR10[4:0], main_swapix2_outR10);
  assign main_swapix2_inR11 = {zll_main_swap2_in[1023:0], 5'hb};
  Main_swapix2  instR79 (main_swapix2_inR11[1028:5], main_swapix2_inR11[4:0], main_swapix2_outR11);
  assign main_swapix2_inR12 = {zll_main_swap2_in[1023:0], 5'hc};
  Main_swapix2  instR80 (main_swapix2_inR12[1028:5], main_swapix2_inR12[4:0], main_swapix2_outR12);
  assign main_swapix2_inR13 = {zll_main_swap2_in[1023:0], 5'hd};
  Main_swapix2  instR81 (main_swapix2_inR13[1028:5], main_swapix2_inR13[4:0], main_swapix2_outR13);
  assign main_swapix2_inR14 = {zll_main_swap2_in[1023:0], 5'he};
  Main_swapix2  instR82 (main_swapix2_inR14[1028:5], main_swapix2_inR14[4:0], main_swapix2_outR14);
  assign main_swapix2_inR15 = {zll_main_swap2_in[1023:0], 5'hf};
  Main_swapix2  instR83 (main_swapix2_inR15[1028:5], main_swapix2_inR15[4:0], main_swapix2_outR15);
  assign main_swapix2_inR16 = {zll_main_swap2_in[1023:0], 5'h10};
  Main_swapix2  instR84 (main_swapix2_inR16[1028:5], main_swapix2_inR16[4:0], main_swapix2_outR16);
  assign main_swapix2_inR17 = {zll_main_swap2_in[1023:0], 5'h11};
  Main_swapix2  instR85 (main_swapix2_inR17[1028:5], main_swapix2_inR17[4:0], main_swapix2_outR17);
  assign main_swapix2_inR18 = {zll_main_swap2_in[1023:0], 5'h12};
  Main_swapix2  instR86 (main_swapix2_inR18[1028:5], main_swapix2_inR18[4:0], main_swapix2_outR18);
  assign main_swapix2_inR19 = {zll_main_swap2_in[1023:0], 5'h13};
  Main_swapix2  instR87 (main_swapix2_inR19[1028:5], main_swapix2_inR19[4:0], main_swapix2_outR19);
  assign main_swapix2_inR20 = {zll_main_swap2_in[1023:0], 5'h14};
  Main_swapix2  instR88 (main_swapix2_inR20[1028:5], main_swapix2_inR20[4:0], main_swapix2_outR20);
  assign main_swapix2_inR21 = {zll_main_swap2_in[1023:0], 5'h15};
  Main_swapix2  instR89 (main_swapix2_inR21[1028:5], main_swapix2_inR21[4:0], main_swapix2_outR21);
  assign main_swapix2_inR22 = {zll_main_swap2_in[1023:0], 5'h16};
  Main_swapix2  instR90 (main_swapix2_inR22[1028:5], main_swapix2_inR22[4:0], main_swapix2_outR22);
  assign main_swapix2_inR23 = {zll_main_swap2_in[1023:0], 5'h17};
  Main_swapix2  instR91 (main_swapix2_inR23[1028:5], main_swapix2_inR23[4:0], main_swapix2_outR23);
  assign main_swapix2_inR24 = {zll_main_swap2_in[1023:0], 5'h18};
  Main_swapix2  instR92 (main_swapix2_inR24[1028:5], main_swapix2_inR24[4:0], main_swapix2_outR24);
  assign main_swapix2_inR25 = {zll_main_swap2_in[1023:0], 5'h19};
  Main_swapix2  instR93 (main_swapix2_inR25[1028:5], main_swapix2_inR25[4:0], main_swapix2_outR25);
  assign main_swapix2_inR26 = {zll_main_swap2_in[1023:0], 5'h1a};
  Main_swapix2  instR94 (main_swapix2_inR26[1028:5], main_swapix2_inR26[4:0], main_swapix2_outR26);
  assign main_swapix2_inR27 = {zll_main_swap2_in[1023:0], 5'h1b};
  Main_swapix2  instR95 (main_swapix2_inR27[1028:5], main_swapix2_inR27[4:0], main_swapix2_outR27);
  assign main_swapix2_inR28 = {zll_main_swap2_in[1023:0], 5'h1c};
  Main_swapix2  instR96 (main_swapix2_inR28[1028:5], main_swapix2_inR28[4:0], main_swapix2_outR28);
  assign main_swapix2_inR29 = {zll_main_swap2_in[1023:0], 5'h1d};
  Main_swapix2  instR97 (main_swapix2_inR29[1028:5], main_swapix2_inR29[4:0], main_swapix2_outR29);
  assign main_swapix2_inR30 = {zll_main_swap2_in[1023:0], 5'h1e};
  Main_swapix2  instR98 (main_swapix2_inR30[1028:5], main_swapix2_inR30[4:0], main_swapix2_outR30);
  assign main_swapix2_inR31 = {zll_main_swap2_in[1023:0], 5'h1f};
  Main_swapix2  instR99 (main_swapix2_inR31[1028:5], main_swapix2_inR31[4:0], main_swapix2_outR31);
  assign zll_main_xor_inR1 = {main_swapix2_out, main_swapix2_outR1, main_swapix2_outR2, main_swapix2_outR3, main_swapix2_outR4, main_swapix2_outR5, main_swapix2_outR6, main_swapix2_outR7, main_swapix2_outR8, main_swapix2_outR9, main_swapix2_outR10, main_swapix2_outR11, main_swapix2_outR12, main_swapix2_outR13, main_swapix2_outR14, main_swapix2_outR15, main_swapix2_outR16, main_swapix2_outR17, main_swapix2_outR18, main_swapix2_outR19, main_swapix2_outR20, main_swapix2_outR21, main_swapix2_outR22, main_swapix2_outR23, main_swapix2_outR24, main_swapix2_outR25, main_swapix2_outR26, main_swapix2_outR27, main_swapix2_outR28, main_swapix2_outR29, main_swapix2_outR30, main_swapix2_outR31};
  ZLL_Main_xor  instR100 (zll_main_xor_inR1[1023:0], zll_main_xor_outR1);
  assign zll_main_swap1_in = zll_main_xor_outR1;
  assign main_swapix1_in = {zll_main_swap1_in[1023:0], 5'h0};
  Main_swapix1  instR101 (main_swapix1_in[1028:5], main_swapix1_in[4:0], main_swapix1_out);
  assign main_swapix1_inR1 = {zll_main_swap1_in[1023:0], 5'h1};
  Main_swapix1  instR102 (main_swapix1_inR1[1028:5], main_swapix1_inR1[4:0], main_swapix1_outR1);
  assign main_swapix1_inR2 = {zll_main_swap1_in[1023:0], 5'h2};
  Main_swapix1  instR103 (main_swapix1_inR2[1028:5], main_swapix1_inR2[4:0], main_swapix1_outR2);
  assign main_swapix1_inR3 = {zll_main_swap1_in[1023:0], 5'h3};
  Main_swapix1  instR104 (main_swapix1_inR3[1028:5], main_swapix1_inR3[4:0], main_swapix1_outR3);
  assign main_swapix1_inR4 = {zll_main_swap1_in[1023:0], 5'h4};
  Main_swapix1  instR105 (main_swapix1_inR4[1028:5], main_swapix1_inR4[4:0], main_swapix1_outR4);
  assign main_swapix1_inR5 = {zll_main_swap1_in[1023:0], 5'h5};
  Main_swapix1  instR106 (main_swapix1_inR5[1028:5], main_swapix1_inR5[4:0], main_swapix1_outR5);
  assign main_swapix1_inR6 = {zll_main_swap1_in[1023:0], 5'h6};
  Main_swapix1  instR107 (main_swapix1_inR6[1028:5], main_swapix1_inR6[4:0], main_swapix1_outR6);
  assign main_swapix1_inR7 = {zll_main_swap1_in[1023:0], 5'h7};
  Main_swapix1  instR108 (main_swapix1_inR7[1028:5], main_swapix1_inR7[4:0], main_swapix1_outR7);
  assign main_swapix1_inR8 = {zll_main_swap1_in[1023:0], 5'h8};
  Main_swapix1  instR109 (main_swapix1_inR8[1028:5], main_swapix1_inR8[4:0], main_swapix1_outR8);
  assign main_swapix1_inR9 = {zll_main_swap1_in[1023:0], 5'h9};
  Main_swapix1  instR110 (main_swapix1_inR9[1028:5], main_swapix1_inR9[4:0], main_swapix1_outR9);
  assign main_swapix1_inR10 = {zll_main_swap1_in[1023:0], 5'ha};
  Main_swapix1  instR111 (main_swapix1_inR10[1028:5], main_swapix1_inR10[4:0], main_swapix1_outR10);
  assign main_swapix1_inR11 = {zll_main_swap1_in[1023:0], 5'hb};
  Main_swapix1  instR112 (main_swapix1_inR11[1028:5], main_swapix1_inR11[4:0], main_swapix1_outR11);
  assign main_swapix1_inR12 = {zll_main_swap1_in[1023:0], 5'hc};
  Main_swapix1  instR113 (main_swapix1_inR12[1028:5], main_swapix1_inR12[4:0], main_swapix1_outR12);
  assign main_swapix1_inR13 = {zll_main_swap1_in[1023:0], 5'hd};
  Main_swapix1  instR114 (main_swapix1_inR13[1028:5], main_swapix1_inR13[4:0], main_swapix1_outR13);
  assign main_swapix1_inR14 = {zll_main_swap1_in[1023:0], 5'he};
  Main_swapix1  instR115 (main_swapix1_inR14[1028:5], main_swapix1_inR14[4:0], main_swapix1_outR14);
  assign main_swapix1_inR15 = {zll_main_swap1_in[1023:0], 5'hf};
  Main_swapix1  instR116 (main_swapix1_inR15[1028:5], main_swapix1_inR15[4:0], main_swapix1_outR15);
  assign main_swapix1_inR16 = {zll_main_swap1_in[1023:0], 5'h10};
  Main_swapix1  instR117 (main_swapix1_inR16[1028:5], main_swapix1_inR16[4:0], main_swapix1_outR16);
  assign main_swapix1_inR17 = {zll_main_swap1_in[1023:0], 5'h11};
  Main_swapix1  instR118 (main_swapix1_inR17[1028:5], main_swapix1_inR17[4:0], main_swapix1_outR17);
  assign main_swapix1_inR18 = {zll_main_swap1_in[1023:0], 5'h12};
  Main_swapix1  instR119 (main_swapix1_inR18[1028:5], main_swapix1_inR18[4:0], main_swapix1_outR18);
  assign main_swapix1_inR19 = {zll_main_swap1_in[1023:0], 5'h13};
  Main_swapix1  instR120 (main_swapix1_inR19[1028:5], main_swapix1_inR19[4:0], main_swapix1_outR19);
  assign main_swapix1_inR20 = {zll_main_swap1_in[1023:0], 5'h14};
  Main_swapix1  instR121 (main_swapix1_inR20[1028:5], main_swapix1_inR20[4:0], main_swapix1_outR20);
  assign main_swapix1_inR21 = {zll_main_swap1_in[1023:0], 5'h15};
  Main_swapix1  instR122 (main_swapix1_inR21[1028:5], main_swapix1_inR21[4:0], main_swapix1_outR21);
  assign main_swapix1_inR22 = {zll_main_swap1_in[1023:0], 5'h16};
  Main_swapix1  instR123 (main_swapix1_inR22[1028:5], main_swapix1_inR22[4:0], main_swapix1_outR22);
  assign main_swapix1_inR23 = {zll_main_swap1_in[1023:0], 5'h17};
  Main_swapix1  instR124 (main_swapix1_inR23[1028:5], main_swapix1_inR23[4:0], main_swapix1_outR23);
  assign main_swapix1_inR24 = {zll_main_swap1_in[1023:0], 5'h18};
  Main_swapix1  instR125 (main_swapix1_inR24[1028:5], main_swapix1_inR24[4:0], main_swapix1_outR24);
  assign main_swapix1_inR25 = {zll_main_swap1_in[1023:0], 5'h19};
  Main_swapix1  instR126 (main_swapix1_inR25[1028:5], main_swapix1_inR25[4:0], main_swapix1_outR25);
  assign main_swapix1_inR26 = {zll_main_swap1_in[1023:0], 5'h1a};
  Main_swapix1  instR127 (main_swapix1_inR26[1028:5], main_swapix1_inR26[4:0], main_swapix1_outR26);
  assign main_swapix1_inR27 = {zll_main_swap1_in[1023:0], 5'h1b};
  Main_swapix1  instR128 (main_swapix1_inR27[1028:5], main_swapix1_inR27[4:0], main_swapix1_outR27);
  assign main_swapix1_inR28 = {zll_main_swap1_in[1023:0], 5'h1c};
  Main_swapix1  instR129 (main_swapix1_inR28[1028:5], main_swapix1_inR28[4:0], main_swapix1_outR28);
  assign main_swapix1_inR29 = {zll_main_swap1_in[1023:0], 5'h1d};
  Main_swapix1  instR130 (main_swapix1_inR29[1028:5], main_swapix1_inR29[4:0], main_swapix1_outR29);
  assign main_swapix1_inR30 = {zll_main_swap1_in[1023:0], 5'h1e};
  Main_swapix1  instR131 (main_swapix1_inR30[1028:5], main_swapix1_inR30[4:0], main_swapix1_outR30);
  assign main_swapix1_inR31 = {zll_main_swap1_in[1023:0], 5'h1f};
  Main_swapix1  instR132 (main_swapix1_inR31[1028:5], main_swapix1_inR31[4:0], main_swapix1_outR31);
  assign main_rotate1_in = {main_swapix1_out, main_swapix1_outR1, main_swapix1_outR2, main_swapix1_outR3, main_swapix1_outR4, main_swapix1_outR5, main_swapix1_outR6, main_swapix1_outR7, main_swapix1_outR8, main_swapix1_outR9, main_swapix1_outR10, main_swapix1_outR11, main_swapix1_outR12, main_swapix1_outR13, main_swapix1_outR14, main_swapix1_outR15, main_swapix1_outR16, main_swapix1_outR17, main_swapix1_outR18, main_swapix1_outR19, main_swapix1_outR20, main_swapix1_outR21, main_swapix1_outR22, main_swapix1_outR23, main_swapix1_outR24, main_swapix1_outR25, main_swapix1_outR26, main_swapix1_outR27, main_swapix1_outR28, main_swapix1_outR29, main_swapix1_outR30, main_swapix1_outR31};
  assign zll_main_rotate_inR1 = {32'h7, main_rotate1_in[1023:0]};
  ZLL_Main_rotate  instR133 (zll_main_rotate_inR1[1055:0], zll_main_rotate_outR1);
  assign zll_main_add_inR1 = zll_main_rotate_outR1;
  ZLL_Main_add  instR134 (zll_main_add_inR1[1023:0], zll_main_add_outR1);
  assign zll_main_nopipeline2_in = zll_main_add_outR1;
  assign zll_main_nopipeline6_in = {{2'h1, {11'h400{1'h0}}}, zll_main_nopipeline2_in[1023:0]};
  assign zll_main_nopipeline24_inR1 = zll_main_nopipeline6_in[2049:0];
  ZLL_Main_nopipeline24  instR135 (zll_main_nopipeline24_inR1[1023:0], zll_main_nopipeline24_outR1);
  assign {__padding, __out0, __st0_next} = (zll_main_nopipeline18_in[0] == 1'h0) ? zll_main_nopipeline24_outR1 : zll_main_nopipeline24_out;
  initial __st0 = {93'h40000000020000001, {10'h3a3{1'h0}}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      __st0 <= {93'h40000000020000001, {10'h3a3{1'h0}}};
    end else begin
      __st0 <= __st0_next;
    end
  end
endmodule

module ZLL_Main_swapix425 (input logic [1023:0] arg0,
  input logic [4:0] arg1,
  output logic [31:0] res);
  logic [4:0] resize_in;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [127:0] resize_inR1;
  logic [2047:0] binop_inR3;
  logic [1023:0] resize_inR2;
  assign resize_in = arg1;
  assign binop_in = {128'h20, 128'(resize_in[4:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h20};
  assign resize_inR1 = binop_inR2[255:128] * binop_inR2[127:0];
  assign binop_inR3 = {arg0, 1024'(resize_inR1[127:0])};
  assign resize_inR2 = binop_inR3[2047:1024] >> binop_inR3[1023:0];
  assign res = resize_inR2[31:0];
endmodule

module Main_rot (input logic [31:0] arg0,
  input logic [1023:0] arg1,
  input logic [4:0] arg2,
  output logic [31:0] res);
  logic [1060:0] zll_main_rot3_in;
  logic [1060:0] zll_main_rot8_in;
  logic [1028:0] main_rotaccess_in;
  logic [1028:0] zll_main_rotaccess3_in;
  logic [1028:0] zll_main_rotaccess12_in;
  logic [4:0] resize_in;
  logic [4:0] zll_main_explode5_in;
  logic [4:0] zll_main_explode5_out;
  logic [1028:0] zll_main_rotaccess1_in;
  logic [1028:0] zll_main_rotaccess10_in;
  logic [1028:0] zll_main_rotaccess5_in;
  logic [1028:0] zll_main_rotaccess9_in;
  logic [4:0] resize_inR1;
  logic [1029:0] zll_main_rotaccess8_in;
  logic [4:0] resize_inR2;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [127:0] resize_inR3;
  logic [2047:0] binop_inR3;
  logic [1023:0] resize_inR4;
  logic [64:0] zll_main_rot10_in;
  logic [64:0] zll_main_rot9_in;
  logic [64:0] zll_main_rot6_in;
  logic [65:0] zll_main_rot2_in;
  logic [64:0] zll_main_rot1_in;
  logic [64:0] zll_main_rot5_in;
  logic [63:0] zll_main_rot12_in;
  logic [63:0] binop_inR4;
  logic [32:0] id_in;
  assign zll_main_rot3_in = {arg0, arg1, arg2};
  assign zll_main_rot8_in = zll_main_rot3_in[1060:0];
  assign main_rotaccess_in = {zll_main_rot8_in[1028:5], zll_main_rot8_in[4:0]};
  assign zll_main_rotaccess3_in = {main_rotaccess_in[1028:5], main_rotaccess_in[4:0]};
  assign zll_main_rotaccess12_in = zll_main_rotaccess3_in[1028:0];
  assign resize_in = zll_main_rotaccess12_in[4:0];
  assign zll_main_explode5_in = resize_in[4:0];
  ZLL_Main_explode5  inst (zll_main_explode5_in[4:0], zll_main_explode5_out);
  assign zll_main_rotaccess1_in = {zll_main_rotaccess12_in[1028:5], zll_main_explode5_out};
  assign zll_main_rotaccess10_in = {zll_main_rotaccess1_in[1028:5], zll_main_rotaccess1_in[4:0]};
  assign zll_main_rotaccess5_in = {zll_main_rotaccess10_in[1028:5], zll_main_rotaccess10_in[3], zll_main_rotaccess10_in[4], zll_main_rotaccess10_in[2], zll_main_rotaccess10_in[1], zll_main_rotaccess10_in[0]};
  assign zll_main_rotaccess9_in = {zll_main_rotaccess5_in[1028:5], zll_main_rotaccess5_in[4], zll_main_rotaccess5_in[3], zll_main_rotaccess5_in[1], zll_main_rotaccess5_in[2], zll_main_rotaccess5_in[0]};
  assign resize_inR1 = {1'h0, zll_main_rotaccess9_in[4], zll_main_rotaccess9_in[1], zll_main_rotaccess9_in[2], zll_main_rotaccess9_in[0]};
  assign zll_main_rotaccess8_in = {zll_main_rotaccess9_in[1028:5], zll_main_rotaccess9_in[3], resize_inR1[4:0]};
  assign resize_inR2 = zll_main_rotaccess8_in[4:0];
  assign binop_in = {128'h20, 128'(resize_inR2[4:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h20};
  assign resize_inR3 = binop_inR2[255:128] * binop_inR2[127:0];
  assign binop_inR3 = {zll_main_rotaccess8_in[1029:6], 1024'(resize_inR3[127:0])};
  assign resize_inR4 = binop_inR3[2047:1024] >> binop_inR3[1023:0];
  assign zll_main_rot10_in = {zll_main_rot8_in[1060:1029], {zll_main_rotaccess8_in[5], resize_inR4[31:0]}};
  assign zll_main_rot9_in = {zll_main_rot10_in[64:33], zll_main_rot10_in[32:0]};
  assign zll_main_rot6_in = {zll_main_rot9_in[32], zll_main_rot9_in[64:33], zll_main_rot9_in[31:0]};
  assign zll_main_rot2_in = {zll_main_rot6_in[64], zll_main_rot6_in[63:32], zll_main_rot6_in[31:0], zll_main_rot6_in[64]};
  assign zll_main_rot1_in = {zll_main_rot2_in[64:33], zll_main_rot2_in[32:1], zll_main_rot2_in[65]};
  assign zll_main_rot5_in = {zll_main_rot1_in[64:33], zll_main_rot1_in[32:1], zll_main_rot1_in[0]};
  assign zll_main_rot12_in = {zll_main_rot5_in[64:33], zll_main_rot5_in[32:1]};
  assign binop_inR4 = {zll_main_rot12_in[31:0], zll_main_rot12_in[63:32]};
  assign id_in = {zll_main_rot2_in[32:1], zll_main_rot2_in[0]};
  assign res = (id_in[0] == 1'h1) ? id_in[32:1] : (binop_inR4[63:32] >>> binop_inR4[31:0]);
endmodule

module ZLL_Main_nopipeline24 (input logic [1023:0] arg0,
  output logic [2049:0] res);
  logic [1023:0] zll_main_nopipeline14_in;
  logic [2047:0] zll_main_nopipeline16_in;
  logic [2047:0] zll_main_nopipeline13_in;
  logic [2049:0] zll_main_nopipeline25_in;
  logic [2049:0] zll_main_nopipeline23_in;
  logic [2047:0] zll_main_nopipeline12_in;
  assign zll_main_nopipeline14_in = arg0;
  assign zll_main_nopipeline16_in = {zll_main_nopipeline14_in[1023:0], zll_main_nopipeline14_in[1023:0]};
  assign zll_main_nopipeline13_in = zll_main_nopipeline16_in[2047:0];
  assign zll_main_nopipeline25_in = {2'h0, zll_main_nopipeline13_in[2047:1024], zll_main_nopipeline13_in[1023:0]};
  assign zll_main_nopipeline23_in = zll_main_nopipeline25_in[2049:0];
  assign zll_main_nopipeline12_in = {zll_main_nopipeline23_in[2047:1024], zll_main_nopipeline23_in[1023:0]};
  assign res = {2'h2, zll_main_nopipeline12_in[2047:1024], zll_main_nopipeline12_in[1023:0]};
endmodule

module ZLL_Main_swapix219 (input logic [4:0] arg0,
  input logic [1023:0] arg1,
  output logic [31:0] res);
  logic [4:0] resize_in;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [127:0] resize_inR1;
  logic [2047:0] binop_inR3;
  logic [1023:0] resize_inR2;
  assign resize_in = arg0;
  assign binop_in = {128'h20, 128'(resize_in[4:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h20};
  assign resize_inR1 = binop_inR2[255:128] * binop_inR2[127:0];
  assign binop_inR3 = {arg1, 1024'(resize_inR1[127:0])};
  assign resize_inR2 = binop_inR3[2047:1024] >> binop_inR3[1023:0];
  assign res = resize_inR2[31:0];
endmodule

module ReWire_Prelude_not (input logic [0:0] arg0,
  output logic [0:0] res);
  logic [1:0] zll_rewire_prelude_not2_in;
  logic [0:0] lit_in;
  assign zll_rewire_prelude_not2_in = {arg0, arg0};
  assign lit_in = zll_rewire_prelude_not2_in[0];
  assign res = (lit_in[0] == 1'h1) ? 1'h0 : 1'h1;
endmodule

module ZLL_Main_add (input logic [1023:0] arg0,
  output logic [1023:0] res);
  logic [1028:0] main_addix_in;
  logic [31:0] main_addix_out;
  logic [1028:0] main_addix_inR1;
  logic [31:0] main_addix_outR1;
  logic [1028:0] main_addix_inR2;
  logic [31:0] main_addix_outR2;
  logic [1028:0] main_addix_inR3;
  logic [31:0] main_addix_outR3;
  logic [1028:0] main_addix_inR4;
  logic [31:0] main_addix_outR4;
  logic [1028:0] main_addix_inR5;
  logic [31:0] main_addix_outR5;
  logic [1028:0] main_addix_inR6;
  logic [31:0] main_addix_outR6;
  logic [1028:0] main_addix_inR7;
  logic [31:0] main_addix_outR7;
  logic [1028:0] main_addix_inR8;
  logic [31:0] main_addix_outR8;
  logic [1028:0] main_addix_inR9;
  logic [31:0] main_addix_outR9;
  logic [1028:0] main_addix_inR10;
  logic [31:0] main_addix_outR10;
  logic [1028:0] main_addix_inR11;
  logic [31:0] main_addix_outR11;
  logic [1028:0] main_addix_inR12;
  logic [31:0] main_addix_outR12;
  logic [1028:0] main_addix_inR13;
  logic [31:0] main_addix_outR13;
  logic [1028:0] main_addix_inR14;
  logic [31:0] main_addix_outR14;
  logic [1028:0] main_addix_inR15;
  logic [31:0] main_addix_outR15;
  logic [1028:0] main_addix_inR16;
  logic [31:0] main_addix_outR16;
  logic [1028:0] main_addix_inR17;
  logic [31:0] main_addix_outR17;
  logic [1028:0] main_addix_inR18;
  logic [31:0] main_addix_outR18;
  logic [1028:0] main_addix_inR19;
  logic [31:0] main_addix_outR19;
  logic [1028:0] main_addix_inR20;
  logic [31:0] main_addix_outR20;
  logic [1028:0] main_addix_inR21;
  logic [31:0] main_addix_outR21;
  logic [1028:0] main_addix_inR22;
  logic [31:0] main_addix_outR22;
  logic [1028:0] main_addix_inR23;
  logic [31:0] main_addix_outR23;
  logic [1028:0] main_addix_inR24;
  logic [31:0] main_addix_outR24;
  logic [1028:0] main_addix_inR25;
  logic [31:0] main_addix_outR25;
  logic [1028:0] main_addix_inR26;
  logic [31:0] main_addix_outR26;
  logic [1028:0] main_addix_inR27;
  logic [31:0] main_addix_outR27;
  logic [1028:0] main_addix_inR28;
  logic [31:0] main_addix_outR28;
  logic [1028:0] main_addix_inR29;
  logic [31:0] main_addix_outR29;
  logic [1028:0] main_addix_inR30;
  logic [31:0] main_addix_outR30;
  logic [1028:0] main_addix_inR31;
  logic [31:0] main_addix_outR31;
  assign main_addix_in = {arg0, 5'h0};
  Main_addix  inst (main_addix_in[1028:5], main_addix_in[4:0], main_addix_out);
  assign main_addix_inR1 = {arg0, 5'h1};
  Main_addix  instR1 (main_addix_inR1[1028:5], main_addix_inR1[4:0], main_addix_outR1);
  assign main_addix_inR2 = {arg0, 5'h2};
  Main_addix  instR2 (main_addix_inR2[1028:5], main_addix_inR2[4:0], main_addix_outR2);
  assign main_addix_inR3 = {arg0, 5'h3};
  Main_addix  instR3 (main_addix_inR3[1028:5], main_addix_inR3[4:0], main_addix_outR3);
  assign main_addix_inR4 = {arg0, 5'h4};
  Main_addix  instR4 (main_addix_inR4[1028:5], main_addix_inR4[4:0], main_addix_outR4);
  assign main_addix_inR5 = {arg0, 5'h5};
  Main_addix  instR5 (main_addix_inR5[1028:5], main_addix_inR5[4:0], main_addix_outR5);
  assign main_addix_inR6 = {arg0, 5'h6};
  Main_addix  instR6 (main_addix_inR6[1028:5], main_addix_inR6[4:0], main_addix_outR6);
  assign main_addix_inR7 = {arg0, 5'h7};
  Main_addix  instR7 (main_addix_inR7[1028:5], main_addix_inR7[4:0], main_addix_outR7);
  assign main_addix_inR8 = {arg0, 5'h8};
  Main_addix  instR8 (main_addix_inR8[1028:5], main_addix_inR8[4:0], main_addix_outR8);
  assign main_addix_inR9 = {arg0, 5'h9};
  Main_addix  instR9 (main_addix_inR9[1028:5], main_addix_inR9[4:0], main_addix_outR9);
  assign main_addix_inR10 = {arg0, 5'ha};
  Main_addix  instR10 (main_addix_inR10[1028:5], main_addix_inR10[4:0], main_addix_outR10);
  assign main_addix_inR11 = {arg0, 5'hb};
  Main_addix  instR11 (main_addix_inR11[1028:5], main_addix_inR11[4:0], main_addix_outR11);
  assign main_addix_inR12 = {arg0, 5'hc};
  Main_addix  instR12 (main_addix_inR12[1028:5], main_addix_inR12[4:0], main_addix_outR12);
  assign main_addix_inR13 = {arg0, 5'hd};
  Main_addix  instR13 (main_addix_inR13[1028:5], main_addix_inR13[4:0], main_addix_outR13);
  assign main_addix_inR14 = {arg0, 5'he};
  Main_addix  instR14 (main_addix_inR14[1028:5], main_addix_inR14[4:0], main_addix_outR14);
  assign main_addix_inR15 = {arg0, 5'hf};
  Main_addix  instR15 (main_addix_inR15[1028:5], main_addix_inR15[4:0], main_addix_outR15);
  assign main_addix_inR16 = {arg0, 5'h10};
  Main_addix  instR16 (main_addix_inR16[1028:5], main_addix_inR16[4:0], main_addix_outR16);
  assign main_addix_inR17 = {arg0, 5'h11};
  Main_addix  instR17 (main_addix_inR17[1028:5], main_addix_inR17[4:0], main_addix_outR17);
  assign main_addix_inR18 = {arg0, 5'h12};
  Main_addix  instR18 (main_addix_inR18[1028:5], main_addix_inR18[4:0], main_addix_outR18);
  assign main_addix_inR19 = {arg0, 5'h13};
  Main_addix  instR19 (main_addix_inR19[1028:5], main_addix_inR19[4:0], main_addix_outR19);
  assign main_addix_inR20 = {arg0, 5'h14};
  Main_addix  instR20 (main_addix_inR20[1028:5], main_addix_inR20[4:0], main_addix_outR20);
  assign main_addix_inR21 = {arg0, 5'h15};
  Main_addix  instR21 (main_addix_inR21[1028:5], main_addix_inR21[4:0], main_addix_outR21);
  assign main_addix_inR22 = {arg0, 5'h16};
  Main_addix  instR22 (main_addix_inR22[1028:5], main_addix_inR22[4:0], main_addix_outR22);
  assign main_addix_inR23 = {arg0, 5'h17};
  Main_addix  instR23 (main_addix_inR23[1028:5], main_addix_inR23[4:0], main_addix_outR23);
  assign main_addix_inR24 = {arg0, 5'h18};
  Main_addix  instR24 (main_addix_inR24[1028:5], main_addix_inR24[4:0], main_addix_outR24);
  assign main_addix_inR25 = {arg0, 5'h19};
  Main_addix  instR25 (main_addix_inR25[1028:5], main_addix_inR25[4:0], main_addix_outR25);
  assign main_addix_inR26 = {arg0, 5'h1a};
  Main_addix  instR26 (main_addix_inR26[1028:5], main_addix_inR26[4:0], main_addix_outR26);
  assign main_addix_inR27 = {arg0, 5'h1b};
  Main_addix  instR27 (main_addix_inR27[1028:5], main_addix_inR27[4:0], main_addix_outR27);
  assign main_addix_inR28 = {arg0, 5'h1c};
  Main_addix  instR28 (main_addix_inR28[1028:5], main_addix_inR28[4:0], main_addix_outR28);
  assign main_addix_inR29 = {arg0, 5'h1d};
  Main_addix  instR29 (main_addix_inR29[1028:5], main_addix_inR29[4:0], main_addix_outR29);
  assign main_addix_inR30 = {arg0, 5'h1e};
  Main_addix  instR30 (main_addix_inR30[1028:5], main_addix_inR30[4:0], main_addix_outR30);
  assign main_addix_inR31 = {arg0, 5'h1f};
  Main_addix  instR31 (main_addix_inR31[1028:5], main_addix_inR31[4:0], main_addix_outR31);
  assign res = {main_addix_out, main_addix_outR1, main_addix_outR2, main_addix_outR3, main_addix_outR4, main_addix_outR5, main_addix_outR6, main_addix_outR7, main_addix_outR8, main_addix_outR9, main_addix_outR10, main_addix_outR11, main_addix_outR12, main_addix_outR13, main_addix_outR14, main_addix_outR15, main_addix_outR16, main_addix_outR17, main_addix_outR18, main_addix_outR19, main_addix_outR20, main_addix_outR21, main_addix_outR22, main_addix_outR23, main_addix_outR24, main_addix_outR25, main_addix_outR26, main_addix_outR27, main_addix_outR28, main_addix_outR29, main_addix_outR30, main_addix_outR31};
endmodule

module Main_swapix4 (input logic [1023:0] arg0,
  input logic [4:0] arg1,
  output logic [31:0] res);
  logic [1028:0] zll_main_swapix47_in;
  logic [1028:0] zll_main_swapix421_in;
  logic [4:0] resize_in;
  logic [4:0] zll_main_explode5_in;
  logic [4:0] zll_main_explode5_out;
  logic [1033:0] zll_main_swapix418_in;
  logic [1033:0] zll_main_swapix423_in;
  logic [1033:0] zll_main_swapix46_in;
  logic [1033:0] zll_main_swapix420_in;
  logic [1033:0] zll_main_swapix424_in;
  logic [4:0] resize_inR1;
  logic [1038:0] zll_main_swapix419_in;
  logic [4:0] resize_inR2;
  logic [1040:0] zll_main_swapix417_in;
  logic [0:0] rewire_prelude_not_in;
  logic [0:0] rewire_prelude_not_out;
  logic [1:0] rewirezupreludezuzazazuin;
  logic [0:0] rewirezupreludezuzaza_out;
  logic [1041:0] zll_main_swapix411_in;
  logic [0:0] rewire_prelude_not_inR1;
  logic [0:0] rewire_prelude_not_outR1;
  logic [1:0] rewirezupreludezuzazazuinR1;
  logic [0:0] rewirezupreludezuzaza_outR1;
  logic [1036:0] zll_main_swapix43_in;
  logic [1036:0] zll_main_swapix48_in;
  logic [1:0] rewirezupreludezuzazazuinR2;
  logic [0:0] rewirezupreludezuzaza_outR2;
  logic [1036:0] zll_main_swapix42_in;
  logic [1:0] rewirezupreludezuzazazuinR3;
  logic [0:0] rewirezupreludezuzaza_outR3;
  logic [1029:0] zll_main_swapix18_in;
  logic [31:0] zll_main_swapix18_out;
  logic [1029:0] zll_main_swapix425_in;
  logic [31:0] zll_main_swapix425_out;
  logic [1029:0] zll_main_swapix425_inR1;
  logic [31:0] zll_main_swapix425_outR1;
  assign zll_main_swapix47_in = {arg0, arg1};
  assign zll_main_swapix421_in = zll_main_swapix47_in[1028:0];
  assign resize_in = zll_main_swapix421_in[4:0];
  assign zll_main_explode5_in = resize_in[4:0];
  ZLL_Main_explode5  inst (zll_main_explode5_in[4:0], zll_main_explode5_out);
  assign zll_main_swapix418_in = {zll_main_swapix421_in[1028:5], zll_main_swapix421_in[4:0], zll_main_explode5_out};
  assign zll_main_swapix423_in = {zll_main_swapix418_in[1033:10], zll_main_swapix418_in[9:5], zll_main_swapix418_in[4:0]};
  assign zll_main_swapix46_in = {zll_main_swapix423_in[4], zll_main_swapix423_in[1033:10], zll_main_swapix423_in[9:5], zll_main_swapix423_in[3], zll_main_swapix423_in[2], zll_main_swapix423_in[1], zll_main_swapix423_in[0]};
  assign zll_main_swapix420_in = {zll_main_swapix46_in[1033], zll_main_swapix46_in[3], zll_main_swapix46_in[1032:9], zll_main_swapix46_in[8:4], zll_main_swapix46_in[2], zll_main_swapix46_in[1], zll_main_swapix46_in[0]};
  assign zll_main_swapix424_in = {zll_main_swapix420_in[1033], zll_main_swapix420_in[1032], zll_main_swapix420_in[1031:8], zll_main_swapix420_in[1], zll_main_swapix420_in[7:3], zll_main_swapix420_in[2], zll_main_swapix420_in[0]};
  assign resize_inR1 = {1'h0, zll_main_swapix424_in[1032], zll_main_swapix424_in[1], zll_main_swapix424_in[7], 1'h1};
  assign zll_main_swapix419_in = {zll_main_swapix424_in[1033], zll_main_swapix424_in[1032], zll_main_swapix424_in[1031:8], zll_main_swapix424_in[0], zll_main_swapix424_in[7], zll_main_swapix424_in[6:2], zll_main_swapix424_in[1], resize_inR1[4:0]};
  assign resize_inR2 = {1'h1, zll_main_swapix419_in[1037], zll_main_swapix419_in[5], zll_main_swapix419_in[11], 1'h0};
  assign zll_main_swapix417_in = {zll_main_swapix419_in[1038], zll_main_swapix419_in[1036:13], zll_main_swapix419_in[12], zll_main_swapix419_in[4:0], zll_main_swapix419_in[10:6], resize_inR2[4:0]};
  assign rewire_prelude_not_in = zll_main_swapix417_in[15];
  ReWire_Prelude_not  instR1 (rewire_prelude_not_in[0], rewire_prelude_not_out);
  assign rewirezupreludezuzazazuin = {zll_main_swapix417_in[1040], rewire_prelude_not_out};
  ReWirezuPreludezuzaza  instR2 (rewirezupreludezuzazazuin[1], rewirezupreludezuzazazuin[0], rewirezupreludezuzaza_out);
  assign zll_main_swapix411_in = {zll_main_swapix417_in[1040], zll_main_swapix417_in[1039:16], zll_main_swapix417_in[15], zll_main_swapix417_in[14:10], zll_main_swapix417_in[9:5], zll_main_swapix417_in[4:0], rewirezupreludezuzaza_out};
  assign rewire_prelude_not_inR1 = zll_main_swapix411_in[16];
  ReWire_Prelude_not  instR3 (rewire_prelude_not_inR1[0], rewire_prelude_not_outR1);
  assign rewirezupreludezuzazazuinR1 = {zll_main_swapix411_in[1041], rewire_prelude_not_outR1};
  ReWirezuPreludezuzaza  instR4 (rewirezupreludezuzazazuinR1[1], rewirezupreludezuzazazuinR1[0], rewirezupreludezuzaza_outR1);
  assign zll_main_swapix43_in = {zll_main_swapix411_in[1041], zll_main_swapix411_in[1040:17], zll_main_swapix411_in[16], zll_main_swapix411_in[10:6], zll_main_swapix411_in[5:1], rewirezupreludezuzaza_outR1};
  assign zll_main_swapix48_in = {zll_main_swapix43_in[1036], zll_main_swapix43_in[1035:12], zll_main_swapix43_in[11], zll_main_swapix43_in[10:6], zll_main_swapix43_in[5:1], zll_main_swapix43_in[0]};
  assign rewirezupreludezuzazazuinR2 = {zll_main_swapix48_in[1036], zll_main_swapix48_in[11]};
  ReWirezuPreludezuzaza  instR5 (rewirezupreludezuzazazuinR2[1], rewirezupreludezuzazazuinR2[0], rewirezupreludezuzaza_outR2);
  assign zll_main_swapix42_in = {zll_main_swapix48_in[1036], zll_main_swapix48_in[1035:12], zll_main_swapix48_in[11], zll_main_swapix48_in[10:6], zll_main_swapix48_in[5:1], rewirezupreludezuzaza_outR2};
  assign rewirezupreludezuzazazuinR3 = {zll_main_swapix42_in[1036], zll_main_swapix42_in[11]};
  ReWirezuPreludezuzaza  instR6 (rewirezupreludezuzazazuinR3[1], rewirezupreludezuzazazuinR3[0], rewirezupreludezuzaza_outR3);
  assign zll_main_swapix18_in = {zll_main_swapix42_in[1035:12], zll_main_swapix42_in[10:6], rewirezupreludezuzaza_outR3};
  ZLL_Main_swapix18  instR7 (zll_main_swapix18_in[1029:6], zll_main_swapix18_in[5:1], zll_main_swapix18_in[0], zll_main_swapix18_out);
  assign zll_main_swapix425_in = {zll_main_swapix42_in[1035:12], zll_main_swapix42_in[5:1], zll_main_swapix42_in[0]};
  ZLL_Main_swapix425  instR8 (zll_main_swapix425_in[1029:6], zll_main_swapix425_in[5:1], zll_main_swapix425_out);
  assign zll_main_swapix425_inR1 = {zll_main_swapix411_in[1040:17], zll_main_swapix411_in[15:11], zll_main_swapix411_in[0]};
  ZLL_Main_swapix425  instR9 (zll_main_swapix425_inR1[1029:6], zll_main_swapix425_inR1[5:1], zll_main_swapix425_outR1);
  assign res = (zll_main_swapix425_inR1[0] == 1'h1) ? zll_main_swapix425_outR1 : ((zll_main_swapix425_in[0] == 1'h1) ? zll_main_swapix425_out : zll_main_swapix18_out);
endmodule

module ZLL_Main_swapix18 (input logic [1023:0] arg0,
  input logic [4:0] arg1,
  input logic [0:0] arg2,
  output logic [31:0] res);
  logic [1029:0] zll_main_swapix416_in;
  logic [1028:0] zll_main_swapix425_in;
  logic [31:0] zll_main_swapix425_out;
  assign zll_main_swapix416_in = {arg0, arg1, arg2};
  assign zll_main_swapix425_in = {zll_main_swapix416_in[1029:6], zll_main_swapix416_in[5:1]};
  ZLL_Main_swapix425  inst (zll_main_swapix425_in[1028:5], zll_main_swapix425_in[4:0], zll_main_swapix425_out);
  assign res = zll_main_swapix425_out;
endmodule

module ZLL_Main_explode5 (input logic [4:0] arg0,
  output logic [4:0] res);
  logic [4:0] resize_in;
  logic [255:0] binop_in;
  logic [127:0] resize_inR1;
  logic [4:0] resize_inR2;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR3;
  logic [4:0] resize_inR4;
  logic [255:0] binop_inR2;
  logic [127:0] resize_inR5;
  logic [4:0] resize_inR6;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR7;
  logic [4:0] resize_inR8;
  logic [255:0] binop_inR4;
  logic [127:0] resize_inR9;
  assign resize_in = arg0;
  assign binop_in = {128'(resize_in[4:0]), 128'h4};
  assign resize_inR1 = binop_in[255:128] >> binop_in[127:0];
  assign resize_inR2 = arg0;
  assign binop_inR1 = {128'(resize_inR2[4:0]), 128'h3};
  assign resize_inR3 = binop_inR1[255:128] >> binop_inR1[127:0];
  assign resize_inR4 = arg0;
  assign binop_inR2 = {128'(resize_inR4[4:0]), 128'h2};
  assign resize_inR5 = binop_inR2[255:128] >> binop_inR2[127:0];
  assign resize_inR6 = arg0;
  assign binop_inR3 = {128'(resize_inR6[4:0]), 128'h1};
  assign resize_inR7 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign resize_inR8 = arg0;
  assign binop_inR4 = {128'(resize_inR8[4:0]), {8'h80{1'h0}}};
  assign resize_inR9 = binop_inR4[255:128] >> binop_inR4[127:0];
  assign res = {resize_inR1[0], resize_inR3[0], resize_inR5[0], resize_inR7[0], resize_inR9[0]};
endmodule

module Main_swapix2 (input logic [1023:0] arg0,
  input logic [4:0] arg1,
  output logic [31:0] res);
  logic [1028:0] zll_main_swapix222_in;
  logic [1028:0] zll_main_swapix210_in;
  logic [4:0] resize_in;
  logic [4:0] zll_main_explode5_in;
  logic [4:0] zll_main_explode5_out;
  logic [1033:0] zll_main_swapix221_in;
  logic [1033:0] zll_main_swapix218_in;
  logic [1033:0] zll_main_swapix2_in;
  logic [1033:0] zll_main_swapix216_in;
  logic [1033:0] zll_main_swapix212_in;
  logic [4:0] resize_inR1;
  logic [1038:0] zll_main_swapix217_in;
  logic [4:0] resize_inR2;
  logic [1040:0] zll_main_swapix215_in;
  logic [0:0] rewire_prelude_not_in;
  logic [0:0] rewire_prelude_not_out;
  logic [1:0] rewirezupreludezuzazazuin;
  logic [0:0] rewirezupreludezuzaza_out;
  logic [1041:0] zll_main_swapix225_in;
  logic [0:0] rewire_prelude_not_inR1;
  logic [0:0] rewire_prelude_not_outR1;
  logic [1:0] rewirezupreludezuzazazuinR1;
  logic [0:0] rewirezupreludezuzaza_outR1;
  logic [1036:0] zll_main_swapix27_in;
  logic [1036:0] zll_main_swapix26_in;
  logic [1:0] rewirezupreludezuzazazuinR2;
  logic [0:0] rewirezupreludezuzaza_outR2;
  logic [1036:0] zll_main_swapix224_in;
  logic [1:0] rewirezupreludezuzazazuinR3;
  logic [0:0] rewirezupreludezuzaza_outR3;
  logic [1029:0] zll_main_swapix24_in;
  logic [1029:0] zll_main_swapix214_in;
  logic [1028:0] zll_main_swapix219_in;
  logic [31:0] zll_main_swapix219_out;
  logic [1029:0] zll_main_swapix219_inR1;
  logic [31:0] zll_main_swapix219_outR1;
  logic [1029:0] zll_main_swapix219_inR2;
  logic [31:0] zll_main_swapix219_outR2;
  assign zll_main_swapix222_in = {arg0, arg1};
  assign zll_main_swapix210_in = zll_main_swapix222_in[1028:0];
  assign resize_in = zll_main_swapix210_in[4:0];
  assign zll_main_explode5_in = resize_in[4:0];
  ZLL_Main_explode5  inst (zll_main_explode5_in[4:0], zll_main_explode5_out);
  assign zll_main_swapix221_in = {zll_main_swapix210_in[4:0], zll_main_swapix210_in[1028:5], zll_main_explode5_out};
  assign zll_main_swapix218_in = {zll_main_swapix221_in[1033:1029], zll_main_swapix221_in[1028:5], zll_main_swapix221_in[4:0]};
  assign zll_main_swapix2_in = {zll_main_swapix218_in[1033:1029], zll_main_swapix218_in[1028:5], zll_main_swapix218_in[3], zll_main_swapix218_in[4], zll_main_swapix218_in[2], zll_main_swapix218_in[1], zll_main_swapix218_in[0]};
  assign zll_main_swapix216_in = {zll_main_swapix2_in[1033:1029], zll_main_swapix2_in[2], zll_main_swapix2_in[1028:5], zll_main_swapix2_in[4], zll_main_swapix2_in[3], zll_main_swapix2_in[1], zll_main_swapix2_in[0]};
  assign zll_main_swapix212_in = {zll_main_swapix216_in[1033:1029], zll_main_swapix216_in[1028], zll_main_swapix216_in[1027:4], zll_main_swapix216_in[3], zll_main_swapix216_in[1], zll_main_swapix216_in[2], zll_main_swapix216_in[0]};
  assign resize_inR1 = {1'h1, zll_main_swapix212_in[3], zll_main_swapix212_in[1028], 1'h1, zll_main_swapix212_in[0]};
  assign zll_main_swapix217_in = {zll_main_swapix212_in[1033:1029], zll_main_swapix212_in[1028], zll_main_swapix212_in[1027:4], zll_main_swapix212_in[3], zll_main_swapix212_in[2], zll_main_swapix212_in[0], zll_main_swapix212_in[1], resize_inR1[4:0]};
  assign resize_inR2 = {1'h1, zll_main_swapix217_in[8], zll_main_swapix217_in[1033], 1'h0, zll_main_swapix217_in[6]};
  assign zll_main_swapix215_in = {zll_main_swapix217_in[4:0], zll_main_swapix217_in[1038:1034], zll_main_swapix217_in[1032:9], zll_main_swapix217_in[7], zll_main_swapix217_in[5], resize_inR2[4:0]};
  assign rewire_prelude_not_in = zll_main_swapix215_in[6];
  ReWire_Prelude_not  instR1 (rewire_prelude_not_in[0], rewire_prelude_not_out);
  assign rewirezupreludezuzazazuin = {zll_main_swapix215_in[5], rewire_prelude_not_out};
  ReWirezuPreludezuzaza  instR2 (rewirezupreludezuzazazuin[1], rewirezupreludezuzazazuin[0], rewirezupreludezuzaza_out);
  assign zll_main_swapix225_in = {zll_main_swapix215_in[1040:1036], zll_main_swapix215_in[4:0], zll_main_swapix215_in[1035:1031], zll_main_swapix215_in[1030:7], zll_main_swapix215_in[6], zll_main_swapix215_in[5], rewirezupreludezuzaza_out};
  assign rewire_prelude_not_inR1 = zll_main_swapix225_in[2];
  ReWire_Prelude_not  instR3 (rewire_prelude_not_inR1[0], rewire_prelude_not_outR1);
  assign rewirezupreludezuzazazuinR1 = {zll_main_swapix225_in[1], rewire_prelude_not_outR1};
  ReWirezuPreludezuzaza  instR4 (rewirezupreludezuzazazuinR1[1], rewirezupreludezuzazazuinR1[0], rewirezupreludezuzaza_outR1);
  assign zll_main_swapix27_in = {zll_main_swapix225_in[1036:1032], zll_main_swapix225_in[1031:1027], zll_main_swapix225_in[1026:3], zll_main_swapix225_in[2], zll_main_swapix225_in[1], rewirezupreludezuzaza_outR1};
  assign zll_main_swapix26_in = {zll_main_swapix27_in[1036:1032], zll_main_swapix27_in[1031:1027], zll_main_swapix27_in[1026:3], zll_main_swapix27_in[2], zll_main_swapix27_in[1], zll_main_swapix27_in[0]};
  assign rewirezupreludezuzazazuinR2 = {zll_main_swapix26_in[1], zll_main_swapix26_in[2]};
  ReWirezuPreludezuzaza  instR5 (rewirezupreludezuzazazuinR2[1], rewirezupreludezuzazazuinR2[0], rewirezupreludezuzaza_outR2);
  assign zll_main_swapix224_in = {zll_main_swapix26_in[1036:1032], zll_main_swapix26_in[1031:1027], zll_main_swapix26_in[1026:3], zll_main_swapix26_in[2], zll_main_swapix26_in[1], rewirezupreludezuzaza_outR2};
  assign rewirezupreludezuzazazuinR3 = {zll_main_swapix224_in[1], zll_main_swapix224_in[2]};
  ReWirezuPreludezuzaza  instR6 (rewirezupreludezuzazazuinR3[1], rewirezupreludezuzazazuinR3[0], rewirezupreludezuzaza_outR3);
  assign zll_main_swapix24_in = {zll_main_swapix224_in[1031:1027], zll_main_swapix224_in[1026:3], rewirezupreludezuzaza_outR3};
  assign zll_main_swapix214_in = {zll_main_swapix24_in[1029:1025], zll_main_swapix24_in[1024:1], zll_main_swapix24_in[0]};
  assign zll_main_swapix219_in = {zll_main_swapix214_in[1029:1025], zll_main_swapix214_in[1024:1]};
  ZLL_Main_swapix219  instR7 (zll_main_swapix219_in[1028:1024], zll_main_swapix219_in[1023:0], zll_main_swapix219_out);
  assign zll_main_swapix219_inR1 = {zll_main_swapix224_in[1036:1032], zll_main_swapix224_in[1026:3], zll_main_swapix224_in[0]};
  ZLL_Main_swapix219  instR8 (zll_main_swapix219_inR1[1029:1025], zll_main_swapix219_inR1[1024:1], zll_main_swapix219_outR1);
  assign zll_main_swapix219_inR2 = {zll_main_swapix225_in[1041:1037], zll_main_swapix225_in[1026:3], zll_main_swapix225_in[0]};
  ZLL_Main_swapix219  instR9 (zll_main_swapix219_inR2[1029:1025], zll_main_swapix219_inR2[1024:1], zll_main_swapix219_outR2);
  assign res = (zll_main_swapix219_inR2[0] == 1'h1) ? zll_main_swapix219_outR2 : ((zll_main_swapix219_inR1[0] == 1'h1) ? zll_main_swapix219_outR1 : zll_main_swapix219_out);
endmodule

module Main_xorix (input logic [1023:0] arg0,
  input logic [4:0] arg1,
  output logic [31:0] res);
  logic [1028:0] zll_main_xorix17_in;
  logic [1028:0] zll_main_xorix6_in;
  logic [4:0] resize_in;
  logic [4:0] zll_main_explode5_in;
  logic [4:0] zll_main_explode5_out;
  logic [1028:0] zll_main_xorix11_in;
  logic [1028:0] zll_main_xorix2_in;
  logic [1028:0] zll_main_xorix1_in;
  logic [1028:0] zll_main_xorix15_in;
  logic [1028:0] zll_main_xorix9_in;
  logic [4:0] resize_inR1;
  logic [1033:0] zll_main_xorix_in;
  logic [4:0] resize_inR2;
  logic [1034:0] zll_main_xorix10_in;
  logic [0:0] rewire_prelude_not_in;
  logic [0:0] rewire_prelude_not_out;
  logic [1035:0] zll_main_xorix7_in;
  logic [0:0] rewire_prelude_not_inR1;
  logic [0:0] rewire_prelude_not_outR1;
  logic [1029:0] zll_main_xorix3_in;
  logic [1029:0] zll_main_swapix425_in;
  logic [31:0] zll_main_swapix425_out;
  logic [1034:0] zll_main_xorix18_in;
  logic [4:0] resize_inR3;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [127:0] resize_inR4;
  logic [2047:0] binop_inR3;
  logic [1023:0] resize_inR5;
  logic [4:0] resize_inR6;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [127:0] resize_inR7;
  logic [2047:0] binop_inR7;
  logic [1023:0] resize_inR8;
  logic [63:0] binop_inR8;
  assign zll_main_xorix17_in = {arg0, arg1};
  assign zll_main_xorix6_in = zll_main_xorix17_in[1028:0];
  assign resize_in = zll_main_xorix6_in[4:0];
  assign zll_main_explode5_in = resize_in[4:0];
  ZLL_Main_explode5  inst (zll_main_explode5_in[4:0], zll_main_explode5_out);
  assign zll_main_xorix11_in = {zll_main_xorix6_in[1028:5], zll_main_explode5_out};
  assign zll_main_xorix2_in = {zll_main_xorix11_in[1028:5], zll_main_xorix11_in[4:0]};
  assign zll_main_xorix1_in = {zll_main_xorix2_in[1028:5], zll_main_xorix2_in[3], zll_main_xorix2_in[4], zll_main_xorix2_in[2], zll_main_xorix2_in[1], zll_main_xorix2_in[0]};
  assign zll_main_xorix15_in = {zll_main_xorix1_in[1028:5], zll_main_xorix1_in[4], zll_main_xorix1_in[2], zll_main_xorix1_in[3], zll_main_xorix1_in[1], zll_main_xorix1_in[0]};
  assign zll_main_xorix9_in = {zll_main_xorix15_in[1028:5], zll_main_xorix15_in[4], zll_main_xorix15_in[1], zll_main_xorix15_in[3], zll_main_xorix15_in[2], zll_main_xorix15_in[0]};
  assign resize_inR1 = {1'h0, zll_main_xorix9_in[4], zll_main_xorix9_in[2], zll_main_xorix9_in[3], zll_main_xorix9_in[0]};
  assign zll_main_xorix_in = {zll_main_xorix9_in[1028:5], zll_main_xorix9_in[4], zll_main_xorix9_in[0], zll_main_xorix9_in[3], zll_main_xorix9_in[2], zll_main_xorix9_in[1], resize_inR1[4:0]};
  assign resize_inR2 = {1'h1, zll_main_xorix_in[9], zll_main_xorix_in[6], zll_main_xorix_in[7], zll_main_xorix_in[8]};
  assign zll_main_xorix10_in = {zll_main_xorix_in[1033:10], zll_main_xorix_in[5], zll_main_xorix_in[4:0], resize_inR2[4:0]};
  assign rewire_prelude_not_in = zll_main_xorix10_in[10];
  ReWire_Prelude_not  instR1 (rewire_prelude_not_in[0], rewire_prelude_not_out);
  assign zll_main_xorix7_in = {zll_main_xorix10_in[1034:11], zll_main_xorix10_in[4:0], zll_main_xorix10_in[10], zll_main_xorix10_in[9:5], rewire_prelude_not_out};
  assign rewire_prelude_not_inR1 = zll_main_xorix7_in[6];
  ReWire_Prelude_not  instR2 (rewire_prelude_not_inR1[0], rewire_prelude_not_outR1);
  assign zll_main_xorix3_in = {zll_main_xorix7_in[1035:12], zll_main_xorix7_in[5:1], rewire_prelude_not_outR1};
  assign zll_main_swapix425_in = {zll_main_xorix3_in[1029:6], zll_main_xorix3_in[5:1], zll_main_xorix3_in[0]};
  ZLL_Main_swapix425  instR3 (zll_main_swapix425_in[1029:6], zll_main_swapix425_in[5:1], zll_main_swapix425_out);
  assign zll_main_xorix18_in = {zll_main_xorix7_in[1035:12], zll_main_xorix7_in[11:7], zll_main_xorix7_in[5:1], zll_main_xorix7_in[0]};
  assign resize_inR3 = zll_main_xorix18_in[5:1];
  assign binop_in = {128'h20, 128'(resize_inR3[4:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h20};
  assign resize_inR4 = binop_inR2[255:128] * binop_inR2[127:0];
  assign binop_inR3 = {zll_main_xorix18_in[1034:11], 1024'(resize_inR4[127:0])};
  assign resize_inR5 = binop_inR3[2047:1024] >> binop_inR3[1023:0];
  assign resize_inR6 = zll_main_xorix18_in[10:6];
  assign binop_inR4 = {128'h20, 128'(resize_inR6[4:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h20};
  assign resize_inR7 = binop_inR6[255:128] * binop_inR6[127:0];
  assign binop_inR7 = {zll_main_xorix18_in[1034:11], 1024'(resize_inR7[127:0])};
  assign resize_inR8 = binop_inR7[2047:1024] >> binop_inR7[1023:0];
  assign binop_inR8 = {resize_inR5[31:0], resize_inR8[31:0]};
  assign res = (zll_main_xorix18_in[0] == 1'h1) ? (binop_inR8[63:32] ^ binop_inR8[31:0]) : zll_main_swapix425_out;
endmodule

module ReWirezuPreludezuzaza (input logic [0:0] arg0,
  input logic [0:0] arg1,
  output logic [0:0] res);
  logic [3:0] zzllzurewirezupreludezuzaza1zuin;
  logic [1:0] zzllzurewirezupreludezuzaza2zuin;
  logic [1:0] lit_in;
  logic [1:0] id_in;
  assign zzllzurewirezupreludezuzaza1zuin = {arg0, arg1, arg0, arg1};
  assign zzllzurewirezupreludezuzaza2zuin = {zzllzurewirezupreludezuzaza1zuin[3], zzllzurewirezupreludezuzaza1zuin[2]};
  assign lit_in = zzllzurewirezupreludezuzaza2zuin[1:0];
  assign id_in = zzllzurewirezupreludezuzaza1zuin[1:0];
  assign res = (id_in[1] == 1'h1) ? id_in[0] : 1'h0;
endmodule

module Main_swapix3 (input logic [1023:0] arg0,
  input logic [4:0] arg1,
  output logic [31:0] res);
  logic [1028:0] zll_main_swapix34_in;
  logic [1028:0] zll_main_swapix321_in;
  logic [4:0] resize_in;
  logic [4:0] zll_main_explode5_in;
  logic [4:0] zll_main_explode5_out;
  logic [1033:0] zll_main_swapix319_in;
  logic [1033:0] zll_main_swapix325_in;
  logic [1033:0] zll_main_swapix320_in;
  logic [1033:0] zll_main_swapix316_in;
  logic [4:0] resize_inR1;
  logic [1038:0] zll_main_swapix314_in;
  logic [4:0] resize_inR2;
  logic [1040:0] zll_main_swapix312_in;
  logic [0:0] rewire_prelude_not_in;
  logic [0:0] rewire_prelude_not_out;
  logic [0:0] rewire_prelude_not_inR1;
  logic [0:0] rewire_prelude_not_outR1;
  logic [1:0] rewirezupreludezuzazazuin;
  logic [0:0] rewirezupreludezuzaza_out;
  logic [1041:0] zll_main_swapix39_in;
  logic [0:0] rewire_prelude_not_inR2;
  logic [0:0] rewire_prelude_not_outR2;
  logic [0:0] rewire_prelude_not_inR3;
  logic [0:0] rewire_prelude_not_outR3;
  logic [1:0] rewirezupreludezuzazazuinR1;
  logic [0:0] rewirezupreludezuzaza_outR1;
  logic [1036:0] zll_main_swapix32_in;
  logic [1036:0] zll_main_swapix33_in;
  logic [0:0] rewire_prelude_not_inR4;
  logic [0:0] rewire_prelude_not_outR4;
  logic [1:0] rewirezupreludezuzazazuinR2;
  logic [0:0] rewirezupreludezuzaza_outR2;
  logic [1036:0] zll_main_swapix322_in;
  logic [0:0] rewire_prelude_not_inR5;
  logic [0:0] rewire_prelude_not_outR5;
  logic [1:0] rewirezupreludezuzazazuinR3;
  logic [0:0] rewirezupreludezuzaza_outR3;
  logic [1029:0] zll_main_swapix18_in;
  logic [31:0] zll_main_swapix18_out;
  logic [1029:0] zll_main_swapix425_in;
  logic [31:0] zll_main_swapix425_out;
  logic [1029:0] zll_main_swapix425_inR1;
  logic [31:0] zll_main_swapix425_outR1;
  assign zll_main_swapix34_in = {arg0, arg1};
  assign zll_main_swapix321_in = zll_main_swapix34_in[1028:0];
  assign resize_in = zll_main_swapix321_in[4:0];
  assign zll_main_explode5_in = resize_in[4:0];
  ZLL_Main_explode5  inst (zll_main_explode5_in[4:0], zll_main_explode5_out);
  assign zll_main_swapix319_in = {zll_main_swapix321_in[1028:5], zll_main_swapix321_in[4:0], zll_main_explode5_out};
  assign zll_main_swapix325_in = {zll_main_swapix319_in[1033:10], zll_main_swapix319_in[9:5], zll_main_swapix319_in[4:0]};
  assign zll_main_swapix320_in = {zll_main_swapix325_in[1033:10], zll_main_swapix325_in[2], zll_main_swapix325_in[9:5], zll_main_swapix325_in[4], zll_main_swapix325_in[3], zll_main_swapix325_in[1], zll_main_swapix325_in[0]};
  assign zll_main_swapix316_in = {zll_main_swapix320_in[1033:10], zll_main_swapix320_in[9], zll_main_swapix320_in[8:4], zll_main_swapix320_in[1], zll_main_swapix320_in[3], zll_main_swapix320_in[2], zll_main_swapix320_in[0]};
  assign resize_inR1 = {1'h0, zll_main_swapix316_in[1], 1'h1, zll_main_swapix316_in[3], zll_main_swapix316_in[0]};
  assign zll_main_swapix314_in = {zll_main_swapix316_in[1033:10], zll_main_swapix316_in[9], zll_main_swapix316_in[0], zll_main_swapix316_in[8:4], zll_main_swapix316_in[3], zll_main_swapix316_in[2], zll_main_swapix316_in[1], resize_inR1[4:0]};
  assign resize_inR2 = {1'h0, zll_main_swapix314_in[5], 1'h0, zll_main_swapix314_in[7], zll_main_swapix314_in[13]};
  assign zll_main_swapix312_in = {zll_main_swapix314_in[1038:15], zll_main_swapix314_in[14], zll_main_swapix314_in[12:8], zll_main_swapix314_in[4:0], zll_main_swapix314_in[6], resize_inR2[4:0]};
  assign rewire_prelude_not_in = zll_main_swapix312_in[5];
  ReWire_Prelude_not  instR1 (rewire_prelude_not_in[0], rewire_prelude_not_out);
  assign rewire_prelude_not_inR1 = zll_main_swapix312_in[16];
  ReWire_Prelude_not  instR2 (rewire_prelude_not_inR1[0], rewire_prelude_not_outR1);
  assign rewirezupreludezuzazazuin = {rewire_prelude_not_out, rewire_prelude_not_outR1};
  ReWirezuPreludezuzaza  instR3 (rewirezupreludezuzazazuin[1], rewirezupreludezuzazazuin[0], rewirezupreludezuzaza_out);
  assign zll_main_swapix39_in = {zll_main_swapix312_in[1040:17], zll_main_swapix312_in[16], zll_main_swapix312_in[15:11], zll_main_swapix312_in[4:0], zll_main_swapix312_in[10:6], zll_main_swapix312_in[5], rewirezupreludezuzaza_out};
  assign rewire_prelude_not_inR2 = zll_main_swapix39_in[1];
  ReWire_Prelude_not  instR4 (rewire_prelude_not_inR2[0], rewire_prelude_not_outR2);
  assign rewire_prelude_not_inR3 = zll_main_swapix39_in[17];
  ReWire_Prelude_not  instR5 (rewire_prelude_not_inR3[0], rewire_prelude_not_outR3);
  assign rewirezupreludezuzazazuinR1 = {rewire_prelude_not_outR2, rewire_prelude_not_outR3};
  ReWirezuPreludezuzaza  instR6 (rewirezupreludezuzazazuinR1[1], rewirezupreludezuzazazuinR1[0], rewirezupreludezuzaza_outR1);
  assign zll_main_swapix32_in = {zll_main_swapix39_in[1041:18], zll_main_swapix39_in[17], zll_main_swapix39_in[16:12], zll_main_swapix39_in[11:7], zll_main_swapix39_in[1], rewirezupreludezuzaza_outR1};
  assign zll_main_swapix33_in = {zll_main_swapix32_in[1036:13], zll_main_swapix32_in[12], zll_main_swapix32_in[11:7], zll_main_swapix32_in[6:2], zll_main_swapix32_in[1], zll_main_swapix32_in[0]};
  assign rewire_prelude_not_inR4 = zll_main_swapix33_in[1];
  ReWire_Prelude_not  instR7 (rewire_prelude_not_inR4[0], rewire_prelude_not_outR4);
  assign rewirezupreludezuzazazuinR2 = {rewire_prelude_not_outR4, zll_main_swapix33_in[12]};
  ReWirezuPreludezuzaza  instR8 (rewirezupreludezuzazazuinR2[1], rewirezupreludezuzazazuinR2[0], rewirezupreludezuzaza_outR2);
  assign zll_main_swapix322_in = {zll_main_swapix33_in[1036:13], zll_main_swapix33_in[12], zll_main_swapix33_in[11:7], zll_main_swapix33_in[6:2], zll_main_swapix33_in[1], rewirezupreludezuzaza_outR2};
  assign rewire_prelude_not_inR5 = zll_main_swapix322_in[1];
  ReWire_Prelude_not  instR9 (rewire_prelude_not_inR5[0], rewire_prelude_not_outR5);
  assign rewirezupreludezuzazazuinR3 = {rewire_prelude_not_outR5, zll_main_swapix322_in[12]};
  ReWirezuPreludezuzaza  instR10 (rewirezupreludezuzazazuinR3[1], rewirezupreludezuzazazuinR3[0], rewirezupreludezuzaza_outR3);
  assign zll_main_swapix18_in = {zll_main_swapix322_in[1036:13], zll_main_swapix322_in[11:7], rewirezupreludezuzaza_outR3};
  ZLL_Main_swapix18  instR11 (zll_main_swapix18_in[1029:6], zll_main_swapix18_in[5:1], zll_main_swapix18_in[0], zll_main_swapix18_out);
  assign zll_main_swapix425_in = {zll_main_swapix322_in[1036:13], zll_main_swapix322_in[6:2], zll_main_swapix322_in[0]};
  ZLL_Main_swapix425  instR12 (zll_main_swapix425_in[1029:6], zll_main_swapix425_in[5:1], zll_main_swapix425_out);
  assign zll_main_swapix425_inR1 = {zll_main_swapix39_in[1041:18], zll_main_swapix39_in[6:2], zll_main_swapix39_in[0]};
  ZLL_Main_swapix425  instR13 (zll_main_swapix425_inR1[1029:6], zll_main_swapix425_inR1[5:1], zll_main_swapix425_outR1);
  assign res = (zll_main_swapix425_inR1[0] == 1'h1) ? zll_main_swapix425_outR1 : ((zll_main_swapix425_in[0] == 1'h1) ? zll_main_swapix425_out : zll_main_swapix18_out);
endmodule

module ZLL_Main_xor (input logic [1023:0] arg0,
  output logic [1023:0] res);
  logic [1028:0] main_xorix_in;
  logic [31:0] main_xorix_out;
  logic [1028:0] main_xorix_inR1;
  logic [31:0] main_xorix_outR1;
  logic [1028:0] main_xorix_inR2;
  logic [31:0] main_xorix_outR2;
  logic [1028:0] main_xorix_inR3;
  logic [31:0] main_xorix_outR3;
  logic [1028:0] main_xorix_inR4;
  logic [31:0] main_xorix_outR4;
  logic [1028:0] main_xorix_inR5;
  logic [31:0] main_xorix_outR5;
  logic [1028:0] main_xorix_inR6;
  logic [31:0] main_xorix_outR6;
  logic [1028:0] main_xorix_inR7;
  logic [31:0] main_xorix_outR7;
  logic [1028:0] main_xorix_inR8;
  logic [31:0] main_xorix_outR8;
  logic [1028:0] main_xorix_inR9;
  logic [31:0] main_xorix_outR9;
  logic [1028:0] main_xorix_inR10;
  logic [31:0] main_xorix_outR10;
  logic [1028:0] main_xorix_inR11;
  logic [31:0] main_xorix_outR11;
  logic [1028:0] main_xorix_inR12;
  logic [31:0] main_xorix_outR12;
  logic [1028:0] main_xorix_inR13;
  logic [31:0] main_xorix_outR13;
  logic [1028:0] main_xorix_inR14;
  logic [31:0] main_xorix_outR14;
  logic [1028:0] main_xorix_inR15;
  logic [31:0] main_xorix_outR15;
  logic [1028:0] main_xorix_inR16;
  logic [31:0] main_xorix_outR16;
  logic [1028:0] main_xorix_inR17;
  logic [31:0] main_xorix_outR17;
  logic [1028:0] main_xorix_inR18;
  logic [31:0] main_xorix_outR18;
  logic [1028:0] main_xorix_inR19;
  logic [31:0] main_xorix_outR19;
  logic [1028:0] main_xorix_inR20;
  logic [31:0] main_xorix_outR20;
  logic [1028:0] main_xorix_inR21;
  logic [31:0] main_xorix_outR21;
  logic [1028:0] main_xorix_inR22;
  logic [31:0] main_xorix_outR22;
  logic [1028:0] main_xorix_inR23;
  logic [31:0] main_xorix_outR23;
  logic [1028:0] main_xorix_inR24;
  logic [31:0] main_xorix_outR24;
  logic [1028:0] main_xorix_inR25;
  logic [31:0] main_xorix_outR25;
  logic [1028:0] main_xorix_inR26;
  logic [31:0] main_xorix_outR26;
  logic [1028:0] main_xorix_inR27;
  logic [31:0] main_xorix_outR27;
  logic [1028:0] main_xorix_inR28;
  logic [31:0] main_xorix_outR28;
  logic [1028:0] main_xorix_inR29;
  logic [31:0] main_xorix_outR29;
  logic [1028:0] main_xorix_inR30;
  logic [31:0] main_xorix_outR30;
  logic [1028:0] main_xorix_inR31;
  logic [31:0] main_xorix_outR31;
  assign main_xorix_in = {arg0, 5'h0};
  Main_xorix  inst (main_xorix_in[1028:5], main_xorix_in[4:0], main_xorix_out);
  assign main_xorix_inR1 = {arg0, 5'h1};
  Main_xorix  instR1 (main_xorix_inR1[1028:5], main_xorix_inR1[4:0], main_xorix_outR1);
  assign main_xorix_inR2 = {arg0, 5'h2};
  Main_xorix  instR2 (main_xorix_inR2[1028:5], main_xorix_inR2[4:0], main_xorix_outR2);
  assign main_xorix_inR3 = {arg0, 5'h3};
  Main_xorix  instR3 (main_xorix_inR3[1028:5], main_xorix_inR3[4:0], main_xorix_outR3);
  assign main_xorix_inR4 = {arg0, 5'h4};
  Main_xorix  instR4 (main_xorix_inR4[1028:5], main_xorix_inR4[4:0], main_xorix_outR4);
  assign main_xorix_inR5 = {arg0, 5'h5};
  Main_xorix  instR5 (main_xorix_inR5[1028:5], main_xorix_inR5[4:0], main_xorix_outR5);
  assign main_xorix_inR6 = {arg0, 5'h6};
  Main_xorix  instR6 (main_xorix_inR6[1028:5], main_xorix_inR6[4:0], main_xorix_outR6);
  assign main_xorix_inR7 = {arg0, 5'h7};
  Main_xorix  instR7 (main_xorix_inR7[1028:5], main_xorix_inR7[4:0], main_xorix_outR7);
  assign main_xorix_inR8 = {arg0, 5'h8};
  Main_xorix  instR8 (main_xorix_inR8[1028:5], main_xorix_inR8[4:0], main_xorix_outR8);
  assign main_xorix_inR9 = {arg0, 5'h9};
  Main_xorix  instR9 (main_xorix_inR9[1028:5], main_xorix_inR9[4:0], main_xorix_outR9);
  assign main_xorix_inR10 = {arg0, 5'ha};
  Main_xorix  instR10 (main_xorix_inR10[1028:5], main_xorix_inR10[4:0], main_xorix_outR10);
  assign main_xorix_inR11 = {arg0, 5'hb};
  Main_xorix  instR11 (main_xorix_inR11[1028:5], main_xorix_inR11[4:0], main_xorix_outR11);
  assign main_xorix_inR12 = {arg0, 5'hc};
  Main_xorix  instR12 (main_xorix_inR12[1028:5], main_xorix_inR12[4:0], main_xorix_outR12);
  assign main_xorix_inR13 = {arg0, 5'hd};
  Main_xorix  instR13 (main_xorix_inR13[1028:5], main_xorix_inR13[4:0], main_xorix_outR13);
  assign main_xorix_inR14 = {arg0, 5'he};
  Main_xorix  instR14 (main_xorix_inR14[1028:5], main_xorix_inR14[4:0], main_xorix_outR14);
  assign main_xorix_inR15 = {arg0, 5'hf};
  Main_xorix  instR15 (main_xorix_inR15[1028:5], main_xorix_inR15[4:0], main_xorix_outR15);
  assign main_xorix_inR16 = {arg0, 5'h10};
  Main_xorix  instR16 (main_xorix_inR16[1028:5], main_xorix_inR16[4:0], main_xorix_outR16);
  assign main_xorix_inR17 = {arg0, 5'h11};
  Main_xorix  instR17 (main_xorix_inR17[1028:5], main_xorix_inR17[4:0], main_xorix_outR17);
  assign main_xorix_inR18 = {arg0, 5'h12};
  Main_xorix  instR18 (main_xorix_inR18[1028:5], main_xorix_inR18[4:0], main_xorix_outR18);
  assign main_xorix_inR19 = {arg0, 5'h13};
  Main_xorix  instR19 (main_xorix_inR19[1028:5], main_xorix_inR19[4:0], main_xorix_outR19);
  assign main_xorix_inR20 = {arg0, 5'h14};
  Main_xorix  instR20 (main_xorix_inR20[1028:5], main_xorix_inR20[4:0], main_xorix_outR20);
  assign main_xorix_inR21 = {arg0, 5'h15};
  Main_xorix  instR21 (main_xorix_inR21[1028:5], main_xorix_inR21[4:0], main_xorix_outR21);
  assign main_xorix_inR22 = {arg0, 5'h16};
  Main_xorix  instR22 (main_xorix_inR22[1028:5], main_xorix_inR22[4:0], main_xorix_outR22);
  assign main_xorix_inR23 = {arg0, 5'h17};
  Main_xorix  instR23 (main_xorix_inR23[1028:5], main_xorix_inR23[4:0], main_xorix_outR23);
  assign main_xorix_inR24 = {arg0, 5'h18};
  Main_xorix  instR24 (main_xorix_inR24[1028:5], main_xorix_inR24[4:0], main_xorix_outR24);
  assign main_xorix_inR25 = {arg0, 5'h19};
  Main_xorix  instR25 (main_xorix_inR25[1028:5], main_xorix_inR25[4:0], main_xorix_outR25);
  assign main_xorix_inR26 = {arg0, 5'h1a};
  Main_xorix  instR26 (main_xorix_inR26[1028:5], main_xorix_inR26[4:0], main_xorix_outR26);
  assign main_xorix_inR27 = {arg0, 5'h1b};
  Main_xorix  instR27 (main_xorix_inR27[1028:5], main_xorix_inR27[4:0], main_xorix_outR27);
  assign main_xorix_inR28 = {arg0, 5'h1c};
  Main_xorix  instR28 (main_xorix_inR28[1028:5], main_xorix_inR28[4:0], main_xorix_outR28);
  assign main_xorix_inR29 = {arg0, 5'h1d};
  Main_xorix  instR29 (main_xorix_inR29[1028:5], main_xorix_inR29[4:0], main_xorix_outR29);
  assign main_xorix_inR30 = {arg0, 5'h1e};
  Main_xorix  instR30 (main_xorix_inR30[1028:5], main_xorix_inR30[4:0], main_xorix_outR30);
  assign main_xorix_inR31 = {arg0, 5'h1f};
  Main_xorix  instR31 (main_xorix_inR31[1028:5], main_xorix_inR31[4:0], main_xorix_outR31);
  assign res = {main_xorix_out, main_xorix_outR1, main_xorix_outR2, main_xorix_outR3, main_xorix_outR4, main_xorix_outR5, main_xorix_outR6, main_xorix_outR7, main_xorix_outR8, main_xorix_outR9, main_xorix_outR10, main_xorix_outR11, main_xorix_outR12, main_xorix_outR13, main_xorix_outR14, main_xorix_outR15, main_xorix_outR16, main_xorix_outR17, main_xorix_outR18, main_xorix_outR19, main_xorix_outR20, main_xorix_outR21, main_xorix_outR22, main_xorix_outR23, main_xorix_outR24, main_xorix_outR25, main_xorix_outR26, main_xorix_outR27, main_xorix_outR28, main_xorix_outR29, main_xorix_outR30, main_xorix_outR31};
endmodule

module Main_swapix1 (input logic [1023:0] arg0,
  input logic [4:0] arg1,
  output logic [31:0] res);
  logic [1028:0] zll_main_swapix16_in;
  logic [1028:0] zll_main_swapix118_in;
  logic [4:0] resize_in;
  logic [4:0] zll_main_explode5_in;
  logic [4:0] zll_main_explode5_out;
  logic [1033:0] zll_main_swapix119_in;
  logic [1033:0] zll_main_swapix121_in;
  logic [1033:0] zll_main_swapix123_in;
  logic [4:0] resize_inR1;
  logic [1038:0] zll_main_swapix120_in;
  logic [4:0] resize_inR2;
  logic [1040:0] zll_main_swapix11_in;
  logic [0:0] rewire_prelude_not_in;
  logic [0:0] rewire_prelude_not_out;
  logic [1:0] rewirezupreludezuzazazuin;
  logic [0:0] rewirezupreludezuzaza_out;
  logic [1041:0] zll_main_swapix115_in;
  logic [0:0] rewire_prelude_not_inR1;
  logic [0:0] rewire_prelude_not_outR1;
  logic [1:0] rewirezupreludezuzazazuinR1;
  logic [0:0] rewirezupreludezuzaza_outR1;
  logic [1036:0] zll_main_swapix111_in;
  logic [1036:0] zll_main_swapix117_in;
  logic [0:0] rewire_prelude_not_inR2;
  logic [0:0] rewire_prelude_not_outR2;
  logic [0:0] rewire_prelude_not_inR3;
  logic [0:0] rewire_prelude_not_outR3;
  logic [1:0] rewirezupreludezuzazazuinR2;
  logic [0:0] rewirezupreludezuzaza_outR2;
  logic [1036:0] zll_main_swapix124_in;
  logic [0:0] rewire_prelude_not_inR4;
  logic [0:0] rewire_prelude_not_outR4;
  logic [0:0] rewire_prelude_not_inR5;
  logic [0:0] rewire_prelude_not_outR5;
  logic [1:0] rewirezupreludezuzazazuinR3;
  logic [0:0] rewirezupreludezuzaza_outR3;
  logic [1029:0] zll_main_swapix18_in;
  logic [31:0] zll_main_swapix18_out;
  logic [1029:0] zll_main_swapix425_in;
  logic [31:0] zll_main_swapix425_out;
  logic [1029:0] zll_main_swapix425_inR1;
  logic [31:0] zll_main_swapix425_outR1;
  assign zll_main_swapix16_in = {arg0, arg1};
  assign zll_main_swapix118_in = zll_main_swapix16_in[1028:0];
  assign resize_in = zll_main_swapix118_in[4:0];
  assign zll_main_explode5_in = resize_in[4:0];
  ZLL_Main_explode5  inst (zll_main_explode5_in[4:0], zll_main_explode5_out);
  assign zll_main_swapix119_in = {zll_main_swapix118_in[1028:5], zll_main_swapix118_in[4:0], zll_main_explode5_out};
  assign zll_main_swapix121_in = {zll_main_swapix119_in[1033:10], zll_main_swapix119_in[9:5], zll_main_swapix119_in[4:0]};
  assign zll_main_swapix123_in = {zll_main_swapix121_in[1033:10], zll_main_swapix121_in[9:5], zll_main_swapix121_in[4], zll_main_swapix121_in[2], zll_main_swapix121_in[3], zll_main_swapix121_in[1], zll_main_swapix121_in[0]};
  assign resize_inR1 = {2'h0, zll_main_swapix123_in[3], zll_main_swapix123_in[1], zll_main_swapix123_in[0]};
  assign zll_main_swapix120_in = {zll_main_swapix123_in[1033:10], zll_main_swapix123_in[9:5], zll_main_swapix123_in[4], zll_main_swapix123_in[3], zll_main_swapix123_in[2], zll_main_swapix123_in[1], zll_main_swapix123_in[0], resize_inR1[4:0]};
  assign resize_inR2 = {2'h1, zll_main_swapix120_in[8], zll_main_swapix120_in[6], zll_main_swapix120_in[5]};
  assign zll_main_swapix11_in = {zll_main_swapix120_in[1038:15], zll_main_swapix120_in[4:0], zll_main_swapix120_in[14:10], zll_main_swapix120_in[9], zll_main_swapix120_in[7], resize_inR2[4:0]};
  assign rewire_prelude_not_in = zll_main_swapix11_in[6];
  ReWire_Prelude_not  instR1 (rewire_prelude_not_in[0], rewire_prelude_not_out);
  assign rewirezupreludezuzazazuin = {rewire_prelude_not_out, zll_main_swapix11_in[5]};
  ReWirezuPreludezuzaza  instR2 (rewirezupreludezuzazazuin[1], rewirezupreludezuzazazuin[0], rewirezupreludezuzaza_out);
  assign zll_main_swapix115_in = {zll_main_swapix11_in[1040:17], zll_main_swapix11_in[16:12], zll_main_swapix11_in[11:7], zll_main_swapix11_in[6], zll_main_swapix11_in[4:0], zll_main_swapix11_in[5], rewirezupreludezuzaza_out};
  assign rewire_prelude_not_inR1 = zll_main_swapix115_in[7];
  ReWire_Prelude_not  instR3 (rewire_prelude_not_inR1[0], rewire_prelude_not_outR1);
  assign rewirezupreludezuzazazuinR1 = {rewire_prelude_not_outR1, zll_main_swapix115_in[1]};
  ReWirezuPreludezuzaza  instR4 (rewirezupreludezuzazazuinR1[1], rewirezupreludezuzazazuinR1[0], rewirezupreludezuzaza_outR1);
  assign zll_main_swapix111_in = {zll_main_swapix115_in[1041:18], zll_main_swapix115_in[12:8], zll_main_swapix115_in[7], zll_main_swapix115_in[6:2], zll_main_swapix115_in[1], rewirezupreludezuzaza_outR1};
  assign zll_main_swapix117_in = {zll_main_swapix111_in[1036:13], zll_main_swapix111_in[12:8], zll_main_swapix111_in[7], zll_main_swapix111_in[6:2], zll_main_swapix111_in[1], zll_main_swapix111_in[0]};
  assign rewire_prelude_not_inR2 = zll_main_swapix117_in[7];
  ReWire_Prelude_not  instR5 (rewire_prelude_not_inR2[0], rewire_prelude_not_outR2);
  assign rewire_prelude_not_inR3 = zll_main_swapix117_in[1];
  ReWire_Prelude_not  instR6 (rewire_prelude_not_inR3[0], rewire_prelude_not_outR3);
  assign rewirezupreludezuzazazuinR2 = {rewire_prelude_not_outR2, rewire_prelude_not_outR3};
  ReWirezuPreludezuzaza  instR7 (rewirezupreludezuzazazuinR2[1], rewirezupreludezuzazazuinR2[0], rewirezupreludezuzaza_outR2);
  assign zll_main_swapix124_in = {zll_main_swapix117_in[1036:13], zll_main_swapix117_in[12:8], zll_main_swapix117_in[7], zll_main_swapix117_in[6:2], zll_main_swapix117_in[1], rewirezupreludezuzaza_outR2};
  assign rewire_prelude_not_inR4 = zll_main_swapix124_in[7];
  ReWire_Prelude_not  instR8 (rewire_prelude_not_inR4[0], rewire_prelude_not_outR4);
  assign rewire_prelude_not_inR5 = zll_main_swapix124_in[1];
  ReWire_Prelude_not  instR9 (rewire_prelude_not_inR5[0], rewire_prelude_not_outR5);
  assign rewirezupreludezuzazazuinR3 = {rewire_prelude_not_outR4, rewire_prelude_not_outR5};
  ReWirezuPreludezuzaza  instR10 (rewirezupreludezuzazazuinR3[1], rewirezupreludezuzazazuinR3[0], rewirezupreludezuzaza_outR3);
  assign zll_main_swapix18_in = {zll_main_swapix124_in[1036:13], zll_main_swapix124_in[12:8], rewirezupreludezuzaza_outR3};
  ZLL_Main_swapix18  instR11 (zll_main_swapix18_in[1029:6], zll_main_swapix18_in[5:1], zll_main_swapix18_in[0], zll_main_swapix18_out);
  assign zll_main_swapix425_in = {zll_main_swapix124_in[1036:13], zll_main_swapix124_in[6:2], zll_main_swapix124_in[0]};
  ZLL_Main_swapix425  instR12 (zll_main_swapix425_in[1029:6], zll_main_swapix425_in[5:1], zll_main_swapix425_out);
  assign zll_main_swapix425_inR1 = {zll_main_swapix115_in[1041:18], zll_main_swapix115_in[17:13], zll_main_swapix115_in[0]};
  ZLL_Main_swapix425  instR13 (zll_main_swapix425_inR1[1029:6], zll_main_swapix425_inR1[5:1], zll_main_swapix425_outR1);
  assign res = (zll_main_swapix425_inR1[0] == 1'h1) ? zll_main_swapix425_outR1 : ((zll_main_swapix425_in[0] == 1'h1) ? zll_main_swapix425_out : zll_main_swapix18_out);
endmodule

module ZLL_Main_rotate (input logic [1055:0] arg0,
  output logic [1023:0] res);
  logic [1055:0] zll_main_rotate2_in;
  logic [1060:0] main_rot_in;
  logic [31:0] main_rot_out;
  logic [1060:0] main_rot_inR1;
  logic [31:0] main_rot_outR1;
  logic [1060:0] main_rot_inR2;
  logic [31:0] main_rot_outR2;
  logic [1060:0] main_rot_inR3;
  logic [31:0] main_rot_outR3;
  logic [1060:0] main_rot_inR4;
  logic [31:0] main_rot_outR4;
  logic [1060:0] main_rot_inR5;
  logic [31:0] main_rot_outR5;
  logic [1060:0] main_rot_inR6;
  logic [31:0] main_rot_outR6;
  logic [1060:0] main_rot_inR7;
  logic [31:0] main_rot_outR7;
  logic [1060:0] main_rot_inR8;
  logic [31:0] main_rot_outR8;
  logic [1060:0] main_rot_inR9;
  logic [31:0] main_rot_outR9;
  logic [1060:0] main_rot_inR10;
  logic [31:0] main_rot_outR10;
  logic [1060:0] main_rot_inR11;
  logic [31:0] main_rot_outR11;
  logic [1060:0] main_rot_inR12;
  logic [31:0] main_rot_outR12;
  logic [1060:0] main_rot_inR13;
  logic [31:0] main_rot_outR13;
  logic [1060:0] main_rot_inR14;
  logic [31:0] main_rot_outR14;
  logic [1060:0] main_rot_inR15;
  logic [31:0] main_rot_outR15;
  logic [1060:0] main_rot_inR16;
  logic [31:0] main_rot_outR16;
  logic [1060:0] main_rot_inR17;
  logic [31:0] main_rot_outR17;
  logic [1060:0] main_rot_inR18;
  logic [31:0] main_rot_outR18;
  logic [1060:0] main_rot_inR19;
  logic [31:0] main_rot_outR19;
  logic [1060:0] main_rot_inR20;
  logic [31:0] main_rot_outR20;
  logic [1060:0] main_rot_inR21;
  logic [31:0] main_rot_outR21;
  logic [1060:0] main_rot_inR22;
  logic [31:0] main_rot_outR22;
  logic [1060:0] main_rot_inR23;
  logic [31:0] main_rot_outR23;
  logic [1060:0] main_rot_inR24;
  logic [31:0] main_rot_outR24;
  logic [1060:0] main_rot_inR25;
  logic [31:0] main_rot_outR25;
  logic [1060:0] main_rot_inR26;
  logic [31:0] main_rot_outR26;
  logic [1060:0] main_rot_inR27;
  logic [31:0] main_rot_outR27;
  logic [1060:0] main_rot_inR28;
  logic [31:0] main_rot_outR28;
  logic [1060:0] main_rot_inR29;
  logic [31:0] main_rot_outR29;
  logic [1060:0] main_rot_inR30;
  logic [31:0] main_rot_outR30;
  logic [1060:0] main_rot_inR31;
  logic [31:0] main_rot_outR31;
  assign zll_main_rotate2_in = arg0;
  assign main_rot_in = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h0};
  Main_rot  inst (main_rot_in[1060:1029], main_rot_in[1028:5], main_rot_in[4:0], main_rot_out);
  assign main_rot_inR1 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h1};
  Main_rot  instR1 (main_rot_inR1[1060:1029], main_rot_inR1[1028:5], main_rot_inR1[4:0], main_rot_outR1);
  assign main_rot_inR2 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h2};
  Main_rot  instR2 (main_rot_inR2[1060:1029], main_rot_inR2[1028:5], main_rot_inR2[4:0], main_rot_outR2);
  assign main_rot_inR3 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h3};
  Main_rot  instR3 (main_rot_inR3[1060:1029], main_rot_inR3[1028:5], main_rot_inR3[4:0], main_rot_outR3);
  assign main_rot_inR4 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h4};
  Main_rot  instR4 (main_rot_inR4[1060:1029], main_rot_inR4[1028:5], main_rot_inR4[4:0], main_rot_outR4);
  assign main_rot_inR5 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h5};
  Main_rot  instR5 (main_rot_inR5[1060:1029], main_rot_inR5[1028:5], main_rot_inR5[4:0], main_rot_outR5);
  assign main_rot_inR6 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h6};
  Main_rot  instR6 (main_rot_inR6[1060:1029], main_rot_inR6[1028:5], main_rot_inR6[4:0], main_rot_outR6);
  assign main_rot_inR7 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h7};
  Main_rot  instR7 (main_rot_inR7[1060:1029], main_rot_inR7[1028:5], main_rot_inR7[4:0], main_rot_outR7);
  assign main_rot_inR8 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h8};
  Main_rot  instR8 (main_rot_inR8[1060:1029], main_rot_inR8[1028:5], main_rot_inR8[4:0], main_rot_outR8);
  assign main_rot_inR9 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h9};
  Main_rot  instR9 (main_rot_inR9[1060:1029], main_rot_inR9[1028:5], main_rot_inR9[4:0], main_rot_outR9);
  assign main_rot_inR10 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'ha};
  Main_rot  instR10 (main_rot_inR10[1060:1029], main_rot_inR10[1028:5], main_rot_inR10[4:0], main_rot_outR10);
  assign main_rot_inR11 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'hb};
  Main_rot  instR11 (main_rot_inR11[1060:1029], main_rot_inR11[1028:5], main_rot_inR11[4:0], main_rot_outR11);
  assign main_rot_inR12 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'hc};
  Main_rot  instR12 (main_rot_inR12[1060:1029], main_rot_inR12[1028:5], main_rot_inR12[4:0], main_rot_outR12);
  assign main_rot_inR13 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'hd};
  Main_rot  instR13 (main_rot_inR13[1060:1029], main_rot_inR13[1028:5], main_rot_inR13[4:0], main_rot_outR13);
  assign main_rot_inR14 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'he};
  Main_rot  instR14 (main_rot_inR14[1060:1029], main_rot_inR14[1028:5], main_rot_inR14[4:0], main_rot_outR14);
  assign main_rot_inR15 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'hf};
  Main_rot  instR15 (main_rot_inR15[1060:1029], main_rot_inR15[1028:5], main_rot_inR15[4:0], main_rot_outR15);
  assign main_rot_inR16 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h10};
  Main_rot  instR16 (main_rot_inR16[1060:1029], main_rot_inR16[1028:5], main_rot_inR16[4:0], main_rot_outR16);
  assign main_rot_inR17 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h11};
  Main_rot  instR17 (main_rot_inR17[1060:1029], main_rot_inR17[1028:5], main_rot_inR17[4:0], main_rot_outR17);
  assign main_rot_inR18 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h12};
  Main_rot  instR18 (main_rot_inR18[1060:1029], main_rot_inR18[1028:5], main_rot_inR18[4:0], main_rot_outR18);
  assign main_rot_inR19 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h13};
  Main_rot  instR19 (main_rot_inR19[1060:1029], main_rot_inR19[1028:5], main_rot_inR19[4:0], main_rot_outR19);
  assign main_rot_inR20 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h14};
  Main_rot  instR20 (main_rot_inR20[1060:1029], main_rot_inR20[1028:5], main_rot_inR20[4:0], main_rot_outR20);
  assign main_rot_inR21 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h15};
  Main_rot  instR21 (main_rot_inR21[1060:1029], main_rot_inR21[1028:5], main_rot_inR21[4:0], main_rot_outR21);
  assign main_rot_inR22 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h16};
  Main_rot  instR22 (main_rot_inR22[1060:1029], main_rot_inR22[1028:5], main_rot_inR22[4:0], main_rot_outR22);
  assign main_rot_inR23 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h17};
  Main_rot  instR23 (main_rot_inR23[1060:1029], main_rot_inR23[1028:5], main_rot_inR23[4:0], main_rot_outR23);
  assign main_rot_inR24 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h18};
  Main_rot  instR24 (main_rot_inR24[1060:1029], main_rot_inR24[1028:5], main_rot_inR24[4:0], main_rot_outR24);
  assign main_rot_inR25 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h19};
  Main_rot  instR25 (main_rot_inR25[1060:1029], main_rot_inR25[1028:5], main_rot_inR25[4:0], main_rot_outR25);
  assign main_rot_inR26 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h1a};
  Main_rot  instR26 (main_rot_inR26[1060:1029], main_rot_inR26[1028:5], main_rot_inR26[4:0], main_rot_outR26);
  assign main_rot_inR27 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h1b};
  Main_rot  instR27 (main_rot_inR27[1060:1029], main_rot_inR27[1028:5], main_rot_inR27[4:0], main_rot_outR27);
  assign main_rot_inR28 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h1c};
  Main_rot  instR28 (main_rot_inR28[1060:1029], main_rot_inR28[1028:5], main_rot_inR28[4:0], main_rot_outR28);
  assign main_rot_inR29 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h1d};
  Main_rot  instR29 (main_rot_inR29[1060:1029], main_rot_inR29[1028:5], main_rot_inR29[4:0], main_rot_outR29);
  assign main_rot_inR30 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h1e};
  Main_rot  instR30 (main_rot_inR30[1060:1029], main_rot_inR30[1028:5], main_rot_inR30[4:0], main_rot_outR30);
  assign main_rot_inR31 = {zll_main_rotate2_in[1055:1024], zll_main_rotate2_in[1023:0], 5'h1f};
  Main_rot  instR31 (main_rot_inR31[1060:1029], main_rot_inR31[1028:5], main_rot_inR31[4:0], main_rot_outR31);
  assign res = {main_rot_out, main_rot_outR1, main_rot_outR2, main_rot_outR3, main_rot_outR4, main_rot_outR5, main_rot_outR6, main_rot_outR7, main_rot_outR8, main_rot_outR9, main_rot_outR10, main_rot_outR11, main_rot_outR12, main_rot_outR13, main_rot_outR14, main_rot_outR15, main_rot_outR16, main_rot_outR17, main_rot_outR18, main_rot_outR19, main_rot_outR20, main_rot_outR21, main_rot_outR22, main_rot_outR23, main_rot_outR24, main_rot_outR25, main_rot_outR26, main_rot_outR27, main_rot_outR28, main_rot_outR29, main_rot_outR30, main_rot_outR31};
endmodule

module Main_addix (input logic [1023:0] arg0,
  input logic [4:0] arg1,
  output logic [31:0] res);
  logic [1028:0] zll_main_addix_in;
  logic [1028:0] zll_main_addix12_in;
  logic [1028:0] main_accesses_in;
  logic [1028:0] zll_main_accesses13_in;
  logic [1028:0] zll_main_accesses4_in;
  logic [4:0] resize_in;
  logic [1028:0] zll_main_accesses2_in;
  logic [4:0] zll_main_explode5_in;
  logic [4:0] zll_main_explode5_out;
  logic [1028:0] zll_main_accesses9_in;
  logic [1028:0] zll_main_accesses1_in;
  logic [1028:0] zll_main_accesses3_in;
  logic [1028:0] zll_main_accesses12_in;
  logic [1028:0] zll_main_accesses8_in;
  logic [4:0] resize_inR1;
  logic [1033:0] zll_main_accesses5_in;
  logic [4:0] resize_inR2;
  logic [1034:0] zll_main_accesses_in;
  logic [4:0] resize_inR3;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [127:0] resize_inR4;
  logic [2047:0] binop_inR3;
  logic [1023:0] resize_inR5;
  logic [4:0] resize_inR6;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [127:0] resize_inR7;
  logic [2047:0] binop_inR7;
  logic [1023:0] resize_inR8;
  logic [64:0] zll_main_addix9_in;
  logic [64:0] zll_main_addix1_in;
  logic [65:0] zll_main_addix6_in;
  logic [32:0] zll_main_addix5_in;
  logic [32:0] id_in;
  logic [64:0] zll_main_addix4_in;
  logic [63:0] binop_inR8;
  assign zll_main_addix_in = {arg0, arg1};
  assign zll_main_addix12_in = zll_main_addix_in[1028:0];
  assign main_accesses_in = {zll_main_addix12_in[1028:5], zll_main_addix12_in[4:0]};
  assign zll_main_accesses13_in = {main_accesses_in[1028:5], main_accesses_in[4:0]};
  assign zll_main_accesses4_in = zll_main_accesses13_in[1028:0];
  assign resize_in = zll_main_accesses4_in[4:0];
  assign zll_main_accesses2_in = {zll_main_accesses4_in[1028:5], resize_in[4:0]};
  assign zll_main_explode5_in = zll_main_accesses2_in[4:0];
  ZLL_Main_explode5  inst (zll_main_explode5_in[4:0], zll_main_explode5_out);
  assign zll_main_accesses9_in = {zll_main_accesses2_in[1028:5], zll_main_explode5_out};
  assign zll_main_accesses1_in = {zll_main_accesses9_in[1028:5], zll_main_accesses9_in[4:0]};
  assign zll_main_accesses3_in = {zll_main_accesses1_in[4], zll_main_accesses1_in[1028:5], zll_main_accesses1_in[3], zll_main_accesses1_in[2], zll_main_accesses1_in[1], zll_main_accesses1_in[0]};
  assign zll_main_accesses12_in = {zll_main_accesses3_in[1028], zll_main_accesses3_in[2], zll_main_accesses3_in[1027:4], zll_main_accesses3_in[3], zll_main_accesses3_in[1], zll_main_accesses3_in[0]};
  assign zll_main_accesses8_in = {zll_main_accesses12_in[1], zll_main_accesses12_in[1028], zll_main_accesses12_in[1027], zll_main_accesses12_in[1026:3], zll_main_accesses12_in[2], zll_main_accesses12_in[0]};
  assign resize_inR1 = {1'h0, zll_main_accesses8_in[1], zll_main_accesses8_in[1026], zll_main_accesses8_in[1028], zll_main_accesses8_in[0]};
  assign zll_main_accesses5_in = {zll_main_accesses8_in[1028], zll_main_accesses8_in[0], zll_main_accesses8_in[1027], zll_main_accesses8_in[1026], zll_main_accesses8_in[1025:2], zll_main_accesses8_in[1], resize_inR1[4:0]};
  assign resize_inR2 = {1'h1, zll_main_accesses5_in[5], zll_main_accesses5_in[1030], zll_main_accesses5_in[1033], zll_main_accesses5_in[1032]};
  assign zll_main_accesses_in = {zll_main_accesses5_in[1031], zll_main_accesses5_in[1029:6], zll_main_accesses5_in[4:0], resize_inR2[4:0]};
  assign resize_inR3 = zll_main_accesses_in[9:5];
  assign binop_in = {128'h20, 128'(resize_inR3[4:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h20};
  assign resize_inR4 = binop_inR2[255:128] * binop_inR2[127:0];
  assign binop_inR3 = {zll_main_accesses_in[1033:10], 1024'(resize_inR4[127:0])};
  assign resize_inR5 = binop_inR3[2047:1024] >> binop_inR3[1023:0];
  assign resize_inR6 = zll_main_accesses_in[4:0];
  assign binop_inR4 = {128'h20, 128'(resize_inR6[4:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h20};
  assign resize_inR7 = binop_inR6[255:128] * binop_inR6[127:0];
  assign binop_inR7 = {zll_main_accesses_in[1033:10], 1024'(resize_inR7[127:0])};
  assign resize_inR8 = binop_inR7[2047:1024] >> binop_inR7[1023:0];
  assign zll_main_addix9_in = {zll_main_accesses_in[1034], resize_inR5[31:0], resize_inR8[31:0]};
  assign zll_main_addix1_in = zll_main_addix9_in[64:0];
  assign zll_main_addix6_in = {zll_main_addix1_in[31:0], zll_main_addix1_in[64], zll_main_addix1_in[63:32], zll_main_addix1_in[64]};
  assign zll_main_addix5_in = {zll_main_addix6_in[32:1], zll_main_addix6_in[33]};
  assign id_in = {zll_main_addix5_in[32:1], zll_main_addix5_in[0]};
  assign zll_main_addix4_in = {zll_main_addix6_in[65:34], zll_main_addix6_in[32:1], zll_main_addix6_in[0]};
  assign binop_inR8 = {zll_main_addix4_in[32:1], zll_main_addix4_in[64:33]};
  assign res = (zll_main_addix4_in[0] == 1'h1) ? (binop_inR8[63:32] + binop_inR8[31:0]) : id_in[32:1];
endmodule