module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [0:0] __in0,
  input logic [31:0] __in1,
  output logic [0:0] __out0,
  output logic [0:0] __out1);
  logic [71:0] zll_pure_dispatch22_in;
  logic [64:0] main_word102_in;
  logic [97:0] zll_main_word1026_in;
  logic [64:0] zll_main_word1023_in;
  logic [64:0] zll_main_word1024_in;
  logic [31:0] zll_main_word1021_in;
  logic [64:0] zll_main_word102_in;
  logic [63:0] zll_main_word1022_in;
  logic [63:0] zll_main_word1025_in;
  logic [71:0] zll_pure_dispatch74_in;
  logic [64:0] main_word24_in;
  logic [97:0] zll_main_word246_in;
  logic [64:0] zll_main_word24_in;
  logic [64:0] zll_main_word245_in;
  logic [31:0] zll_main_word244_in;
  logic [64:0] zll_main_word241_in;
  logic [63:0] zll_main_word242_in;
  logic [63:0] zll_main_word243_in;
  logic [71:0] zll_pure_dispatch20_in;
  logic [64:0] main_word111_in;
  logic [97:0] zll_main_word1115_in;
  logic [64:0] zll_main_word1113_in;
  logic [64:0] zll_main_word111_in;
  logic [31:0] zll_main_word1119_in;
  logic [64:0] zll_main_word1118_in;
  logic [63:0] zll_main_word1112_in;
  logic [63:0] zll_main_word1111_in;
  logic [71:0] zll_pure_dispatch94_in;
  logic [64:0] main_word10_in;
  logic [97:0] zll_main_word1018_in;
  logic [64:0] zll_main_word108_in;
  logic [64:0] zll_main_word1010_in;
  logic [31:0] zll_main_word10_in;
  logic [64:0] zll_main_word1015_in;
  logic [63:0] zll_main_word101_in;
  logic [63:0] zll_main_word1017_in;
  logic [71:0] zll_pure_dispatch5_in;
  logic [64:0] main_word51_in;
  logic [97:0] zll_main_word511_in;
  logic [64:0] zll_main_word518_in;
  logic [64:0] zll_main_word516_in;
  logic [31:0] zll_main_word5111_in;
  logic [64:0] zll_main_word5110_in;
  logic [63:0] zll_main_word512_in;
  logic [63:0] zll_main_word51_in;
  logic [71:0] zll_pure_dispatch45_in;
  logic [64:0] main_word4_in;
  logic [97:0] zll_main_word420_in;
  logic [64:0] zll_main_word41_in;
  logic [64:0] zll_main_word425_in;
  logic [31:0] zll_main_word4_in;
  logic [64:0] zll_main_word423_in;
  logic [63:0] zll_main_word410_in;
  logic [63:0] zll_main_word417_in;
  logic [63:0] zll_main_word430_in;
  logic [65:0] zll_main_word430_out;
  logic [97:0] zll_main_word43_in;
  logic [97:0] zll_main_word428_in;
  logic [95:0] zll_main_word418_in;
  logic [63:0] test2_in;
  logic [0:0] extres;
  logic [71:0] zll_pure_dispatch68_in;
  logic [64:0] main_word71_in;
  logic [97:0] zll_main_word713_in;
  logic [64:0] zll_main_word716_in;
  logic [64:0] zll_main_word712_in;
  logic [31:0] zll_main_word71_in;
  logic [64:0] zll_main_word718_in;
  logic [63:0] zll_main_word711_in;
  logic [63:0] zll_main_word719_in;
  logic [71:0] zll_pure_dispatch123_in;
  logic [64:0] main_word103_in;
  logic [97:0] zll_main_word1036_in;
  logic [64:0] zll_main_word103_in;
  logic [64:0] zll_main_word1031_in;
  logic [31:0] zll_main_word1034_in;
  logic [64:0] zll_main_word1035_in;
  logic [63:0] zll_main_word1033_in;
  logic [63:0] zll_main_word1032_in;
  logic [71:0] zll_pure_dispatch9_in;
  logic [64:0] main_word122_in;
  logic [97:0] zll_main_word1222_in;
  logic [64:0] zll_main_word1226_in;
  logic [64:0] zll_main_word1225_in;
  logic [31:0] zll_main_word1223_in;
  logic [64:0] zll_main_word1224_in;
  logic [63:0] zll_main_word1221_in;
  logic [63:0] zll_main_word122_in;
  logic [71:0] zll_pure_dispatch12_in;
  logic [64:0] main_word126_in;
  logic [97:0] zll_main_word1265_in;
  logic [64:0] zll_main_word126_in;
  logic [64:0] zll_main_word1262_in;
  logic [31:0] zll_main_word1264_in;
  logic [64:0] zll_main_word1263_in;
  logic [63:0] zll_main_word1261_in;
  logic [63:0] zll_main_word1266_in;
  logic [71:0] zll_pure_dispatch124_in;
  logic [64:0] main_word81_in;
  logic [97:0] zll_main_word813_in;
  logic [64:0] zll_main_word818_in;
  logic [64:0] zll_main_word812_in;
  logic [31:0] zll_main_word816_in;
  logic [64:0] zll_main_word811_in;
  logic [63:0] zll_main_word814_in;
  logic [63:0] zll_main_word817_in;
  logic [71:0] zll_pure_dispatch85_in;
  logic [64:0] main_word107_in;
  logic [97:0] zll_main_word1073_in;
  logic [64:0] zll_main_word107_in;
  logic [64:0] zll_main_word1075_in;
  logic [31:0] zll_main_word1071_in;
  logic [64:0] zll_main_word1076_in;
  logic [63:0] zll_main_word1072_in;
  logic [63:0] zll_main_word1074_in;
  logic [71:0] zll_pure_dispatch49_in;
  logic [64:0] main_word118_in;
  logic [97:0] zll_main_word1184_in;
  logic [64:0] zll_main_word1182_in;
  logic [64:0] zll_main_word1187_in;
  logic [31:0] zll_main_word1183_in;
  logic [64:0] zll_main_word1181_in;
  logic [63:0] zll_main_word1185_in;
  logic [63:0] zll_main_word1186_in;
  logic [71:0] zll_pure_dispatch76_in;
  logic [64:0] main_word61_in;
  logic [97:0] zll_main_word616_in;
  logic [64:0] zll_main_word6110_in;
  logic [64:0] zll_main_word612_in;
  logic [31:0] zll_main_word61_in;
  logic [64:0] zll_main_word6112_in;
  logic [63:0] zll_main_word618_in;
  logic [63:0] zll_main_word6111_in;
  logic [71:0] zll_pure_dispatch114_in;
  logic [64:0] main_word98_in;
  logic [97:0] zll_main_word985_in;
  logic [64:0] zll_main_word983_in;
  logic [64:0] zll_main_word986_in;
  logic [31:0] zll_main_word98_in;
  logic [64:0] zll_main_word982_in;
  logic [63:0] zll_main_word981_in;
  logic [63:0] zll_main_word984_in;
  logic [71:0] zll_pure_dispatch10_in;
  logic [64:0] main_word18_in;
  logic [97:0] zll_main_word183_in;
  logic [64:0] zll_main_word185_in;
  logic [64:0] zll_main_word182_in;
  logic [31:0] zll_main_word18_in;
  logic [64:0] zll_main_word186_in;
  logic [63:0] zll_main_word184_in;
  logic [63:0] zll_main_word181_in;
  logic [71:0] zll_pure_dispatch42_in;
  logic [64:0] main_word100_in;
  logic [97:0] zll_main_word1005_in;
  logic [64:0] zll_main_word1004_in;
  logic [64:0] zll_main_word100_in;
  logic [31:0] zll_main_word1006_in;
  logic [64:0] zll_main_word1003_in;
  logic [63:0] zll_main_word1002_in;
  logic [63:0] zll_main_word1001_in;
  logic [71:0] zll_pure_dispatch37_in;
  logic [64:0] main_word125_in;
  logic [97:0] zll_main_word1254_in;
  logic [64:0] zll_main_word1255_in;
  logic [64:0] zll_main_word1252_in;
  logic [31:0] zll_main_word1251_in;
  logic [64:0] zll_main_word1256_in;
  logic [63:0] zll_main_word125_in;
  logic [63:0] zll_main_word1253_in;
  logic [71:0] zll_pure_dispatch96_in;
  logic [64:0] main_word59_in;
  logic [97:0] zll_main_word592_in;
  logic [64:0] zll_main_word596_in;
  logic [64:0] zll_main_word595_in;
  logic [31:0] zll_main_word593_in;
  logic [64:0] zll_main_word594_in;
  logic [63:0] zll_main_word597_in;
  logic [63:0] zll_main_word591_in;
  logic [71:0] zll_pure_dispatch99_in;
  logic [64:0] main_word32_in;
  logic [97:0] zll_main_word327_in;
  logic [64:0] zll_main_word324_in;
  logic [64:0] zll_main_word32_in;
  logic [31:0] zll_main_word322_in;
  logic [64:0] zll_main_word323_in;
  logic [63:0] zll_main_word321_in;
  logic [63:0] zll_main_word325_in;
  logic [71:0] zll_pure_dispatch110_in;
  logic [64:0] main_word68_in;
  logic [97:0] zll_main_word685_in;
  logic [64:0] zll_main_word683_in;
  logic [64:0] zll_main_word682_in;
  logic [31:0] zll_main_word68_in;
  logic [64:0] zll_main_word681_in;
  logic [63:0] zll_main_word684_in;
  logic [63:0] zll_main_word686_in;
  logic [71:0] zll_pure_dispatch93_in;
  logic [64:0] main_word37_in;
  logic [97:0] zll_main_word373_in;
  logic [64:0] zll_main_word377_in;
  logic [64:0] zll_main_word372_in;
  logic [31:0] zll_main_word375_in;
  logic [64:0] zll_main_word374_in;
  logic [63:0] zll_main_word376_in;
  logic [63:0] zll_main_word371_in;
  logic [71:0] zll_pure_dispatch58_in;
  logic [64:0] main_word58_in;
  logic [97:0] zll_main_word586_in;
  logic [64:0] zll_main_word583_in;
  logic [64:0] zll_main_word584_in;
  logic [31:0] zll_main_word58_in;
  logic [64:0] zll_main_word582_in;
  logic [63:0] zll_main_word581_in;
  logic [63:0] zll_main_word585_in;
  logic [71:0] zll_pure_dispatch92_in;
  logic [64:0] main_word31_in;
  logic [97:0] zll_main_word315_in;
  logic [64:0] zll_main_word311_in;
  logic [64:0] zll_main_word3110_in;
  logic [31:0] zll_main_word319_in;
  logic [64:0] zll_main_word31_in;
  logic [63:0] zll_main_word312_in;
  logic [63:0] zll_main_word3111_in;
  logic [71:0] zll_pure_dispatch15_in;
  logic [64:0] main_word82_in;
  logic [97:0] zll_main_word821_in;
  logic [64:0] zll_main_word823_in;
  logic [64:0] zll_main_word824_in;
  logic [31:0] zll_main_word825_in;
  logic [64:0] zll_main_word822_in;
  logic [63:0] zll_main_word826_in;
  logic [63:0] zll_main_word827_in;
  logic [71:0] zll_pure_dispatch86_in;
  logic [64:0] main_word52_in;
  logic [97:0] zll_main_word525_in;
  logic [64:0] zll_main_word524_in;
  logic [64:0] zll_main_word5210_in;
  logic [31:0] zll_main_word521_in;
  logic [64:0] zll_main_word526_in;
  logic [63:0] zll_main_word522_in;
  logic [63:0] zll_main_word523_in;
  logic [71:0] zll_pure_dispatch8_in;
  logic [64:0] main_word101_in;
  logic [97:0] zll_main_word1011_in;
  logic [64:0] zll_main_word1016_in;
  logic [64:0] zll_main_word1019_in;
  logic [31:0] zll_main_word1012_in;
  logic [64:0] zll_main_word10110_in;
  logic [63:0] zll_main_word1014_in;
  logic [63:0] zll_main_word1013_in;
  logic [71:0] zll_pure_dispatch116_in;
  logic [64:0] main_word80_in;
  logic [97:0] zll_main_word803_in;
  logic [64:0] zll_main_word802_in;
  logic [64:0] zll_main_word804_in;
  logic [31:0] zll_main_word801_in;
  logic [64:0] zll_main_word806_in;
  logic [63:0] zll_main_word80_in;
  logic [63:0] zll_main_word805_in;
  logic [71:0] zll_pure_dispatch90_in;
  logic [64:0] main_word39_in;
  logic [97:0] zll_main_word39_in;
  logic [64:0] zll_main_word395_in;
  logic [64:0] zll_main_word393_in;
  logic [31:0] zll_main_word391_in;
  logic [64:0] zll_main_word392_in;
  logic [63:0] zll_main_word394_in;
  logic [63:0] zll_main_word396_in;
  logic [71:0] zll_pure_dispatch7_in;
  logic [64:0] main_word21_in;
  logic [97:0] zll_main_word216_in;
  logic [64:0] zll_main_word2110_in;
  logic [64:0] zll_main_word2112_in;
  logic [31:0] zll_main_word218_in;
  logic [64:0] zll_main_word2111_in;
  logic [63:0] zll_main_word217_in;
  logic [63:0] zll_main_word2113_in;
  logic [71:0] zll_pure_dispatch88_in;
  logic [64:0] main_word16_in;
  logic [97:0] zll_main_word164_in;
  logic [64:0] zll_main_word163_in;
  logic [64:0] zll_main_word162_in;
  logic [31:0] zll_main_word165_in;
  logic [64:0] zll_main_word161_in;
  logic [63:0] zll_main_word166_in;
  logic [63:0] zll_main_word16_in;
  logic [71:0] zll_pure_dispatch97_in;
  logic [64:0] main_word112_in;
  logic [97:0] zll_main_word112_in;
  logic [64:0] zll_main_word1121_in;
  logic [64:0] zll_main_word1123_in;
  logic [31:0] zll_main_word1126_in;
  logic [64:0] zll_main_word1122_in;
  logic [63:0] zll_main_word1124_in;
  logic [63:0] zll_main_word1125_in;
  logic [71:0] zll_pure_dispatch80_in;
  logic [64:0] main_word12_in;
  logic [97:0] zll_main_word124_in;
  logic [64:0] zll_main_word1215_in;
  logic [64:0] zll_main_word1219_in;
  logic [31:0] zll_main_word1210_in;
  logic [64:0] zll_main_word127_in;
  logic [63:0] zll_main_word1211_in;
  logic [63:0] zll_main_word1213_in;
  logic [71:0] zll_pure_dispatch87_in;
  logic [64:0] main_word42_in;
  logic [97:0] zll_main_word429_in;
  logic [64:0] zll_main_word421_in;
  logic [64:0] zll_main_word4210_in;
  logic [31:0] zll_main_word4212_in;
  logic [64:0] zll_main_word42_in;
  logic [63:0] zll_main_word4211_in;
  logic [63:0] zll_main_word424_in;
  logic [71:0] zll_pure_dispatch57_in;
  logic [64:0] main_word1_in;
  logic [97:0] zll_main_word121_in;
  logic [64:0] zll_main_word147_in;
  logic [64:0] zll_main_word09_in;
  logic [65:0] zll_main_word09_out;
  logic [64:0] zll_main_word130_in;
  logic [63:0] zll_main_word138_in;
  logic [63:0] zll_main_word133_in;
  logic [63:0] zll_main_word430_inR1;
  logic [65:0] zll_main_word430_outR1;
  logic [97:0] zll_main_word12_in;
  logic [97:0] zll_main_word140_in;
  logic [95:0] zll_main_word128_in;
  logic [63:0] test1_in;
  logic [0:0] extresR1;
  logic [71:0] zll_pure_dispatch111_in;
  logic [64:0] main_word41_in;
  logic [97:0] zll_main_word413_in;
  logic [64:0] zll_main_word411_in;
  logic [64:0] zll_main_word415_in;
  logic [31:0] zll_main_word416_in;
  logic [64:0] zll_main_word414_in;
  logic [63:0] zll_main_word4110_in;
  logic [63:0] zll_main_word412_in;
  logic [71:0] zll_pure_dispatch32_in;
  logic [64:0] main_word96_in;
  logic [97:0] zll_main_word966_in;
  logic [64:0] zll_main_word961_in;
  logic [64:0] zll_main_word964_in;
  logic [31:0] zll_main_word963_in;
  logic [64:0] zll_main_word965_in;
  logic [63:0] zll_main_word96_in;
  logic [63:0] zll_main_word962_in;
  logic [71:0] zll_pure_dispatch79_in;
  logic [64:0] main_word53_in;
  logic [97:0] zll_main_word535_in;
  logic [64:0] zll_main_word53_in;
  logic [64:0] zll_main_word532_in;
  logic [31:0] zll_main_word533_in;
  logic [64:0] zll_main_word531_in;
  logic [63:0] zll_main_word536_in;
  logic [63:0] zll_main_word534_in;
  logic [71:0] zll_pure_dispatch44_in;
  logic [64:0] main_word89_in;
  logic [97:0] zll_main_word894_in;
  logic [64:0] zll_main_word896_in;
  logic [64:0] zll_main_word892_in;
  logic [31:0] zll_main_word895_in;
  logic [64:0] zll_main_word891_in;
  logic [63:0] zll_main_word89_in;
  logic [63:0] zll_main_word893_in;
  logic [71:0] zll_pure_dispatch82_in;
  logic [64:0] main_word35_in;
  logic [97:0] zll_main_word353_in;
  logic [64:0] zll_main_word35_in;
  logic [64:0] zll_main_word351_in;
  logic [31:0] zll_main_word354_in;
  logic [64:0] zll_main_word352_in;
  logic [63:0] zll_main_word355_in;
  logic [63:0] zll_main_word356_in;
  logic [71:0] zll_pure_dispatch19_in;
  logic [64:0] main_word94_in;
  logic [97:0] zll_main_word94_in;
  logic [64:0] zll_main_word945_in;
  logic [64:0] zll_main_word944_in;
  logic [31:0] zll_main_word946_in;
  logic [64:0] zll_main_word943_in;
  logic [63:0] zll_main_word942_in;
  logic [63:0] zll_main_word941_in;
  logic [71:0] zll_pure_dispatch71_in;
  logic [64:0] main_word55_in;
  logic [97:0] zll_main_word55_in;
  logic [64:0] zll_main_word552_in;
  logic [64:0] zll_main_word551_in;
  logic [31:0] zll_main_word556_in;
  logic [64:0] zll_main_word553_in;
  logic [63:0] zll_main_word555_in;
  logic [63:0] zll_main_word554_in;
  logic [71:0] zll_pure_dispatch48_in;
  logic [64:0] main_word26_in;
  logic [97:0] zll_main_word266_in;
  logic [64:0] zll_main_word264_in;
  logic [64:0] zll_main_word263_in;
  logic [31:0] zll_main_word261_in;
  logic [64:0] zll_main_word26_in;
  logic [63:0] zll_main_word265_in;
  logic [63:0] zll_main_word262_in;
  logic [71:0] zll_pure_dispatch77_in;
  logic [64:0] main_word123_in;
  logic [97:0] zll_main_word1236_in;
  logic [64:0] zll_main_word1231_in;
  logic [64:0] zll_main_word1233_in;
  logic [31:0] zll_main_word1235_in;
  logic [64:0] zll_main_word1232_in;
  logic [63:0] zll_main_word123_in;
  logic [63:0] zll_main_word1234_in;
  logic [71:0] zll_pure_dispatch27_in;
  logic [64:0] main_word27_in;
  logic [97:0] zll_main_word271_in;
  logic [64:0] zll_main_word272_in;
  logic [64:0] zll_main_word27_in;
  logic [31:0] zll_main_word273_in;
  logic [64:0] zll_main_word275_in;
  logic [63:0] zll_main_word274_in;
  logic [63:0] zll_main_word276_in;
  logic [71:0] zll_pure_dispatch41_in;
  logic [64:0] main_word83_in;
  logic [97:0] zll_main_word831_in;
  logic [64:0] zll_main_word835_in;
  logic [64:0] zll_main_word83_in;
  logic [31:0] zll_main_word833_in;
  logic [64:0] zll_main_word836_in;
  logic [63:0] zll_main_word832_in;
  logic [63:0] zll_main_word834_in;
  logic [71:0] zll_pure_dispatch117_in;
  logic [64:0] main_word13_in;
  logic [97:0] zll_main_word137_in;
  logic [64:0] zll_main_word132_in;
  logic [64:0] zll_main_word131_in;
  logic [31:0] zll_main_word134_in;
  logic [64:0] zll_main_word13_in;
  logic [63:0] zll_main_word1311_in;
  logic [63:0] zll_main_word1310_in;
  logic [71:0] zll_pure_dispatch64_in;
  logic [64:0] main_word69_in;
  logic [97:0] zll_main_word695_in;
  logic [64:0] zll_main_word69_in;
  logic [64:0] zll_main_word691_in;
  logic [31:0] zll_main_word693_in;
  logic [64:0] zll_main_word692_in;
  logic [63:0] zll_main_word696_in;
  logic [63:0] zll_main_word694_in;
  logic [71:0] zll_pure_dispatch69_in;
  logic [64:0] main_word115_in;
  logic [97:0] zll_main_word1155_in;
  logic [64:0] zll_main_word1152_in;
  logic [64:0] zll_main_word1153_in;
  logic [31:0] zll_main_word1154_in;
  logic [64:0] zll_main_word1151_in;
  logic [63:0] zll_main_word115_in;
  logic [63:0] zll_main_word1156_in;
  logic [71:0] zll_pure_dispatch21_in;
  logic [64:0] main_word87_in;
  logic [97:0] zll_main_word875_in;
  logic [64:0] zll_main_word873_in;
  logic [64:0] zll_main_word87_in;
  logic [31:0] zll_main_word874_in;
  logic [64:0] zll_main_word872_in;
  logic [63:0] zll_main_word871_in;
  logic [63:0] zll_main_word876_in;
  logic [71:0] zll_pure_dispatch72_in;
  logic [64:0] main_word25_in;
  logic [97:0] zll_main_word254_in;
  logic [64:0] zll_main_word256_in;
  logic [64:0] zll_main_word251_in;
  logic [31:0] zll_main_word252_in;
  logic [64:0] zll_main_word25_in;
  logic [63:0] zll_main_word253_in;
  logic [63:0] zll_main_word255_in;
  logic [71:0] zll_pure_dispatch103_in;
  logic [64:0] main_word19_in;
  logic [97:0] zll_main_word196_in;
  logic [64:0] zll_main_word194_in;
  logic [64:0] zll_main_word193_in;
  logic [31:0] zll_main_word19_in;
  logic [64:0] zll_main_word195_in;
  logic [63:0] zll_main_word191_in;
  logic [63:0] zll_main_word192_in;
  logic [71:0] zll_pure_dispatch62_in;
  logic [64:0] main_word76_in;
  logic [97:0] zll_main_word762_in;
  logic [64:0] zll_main_word765_in;
  logic [64:0] zll_main_word761_in;
  logic [31:0] zll_main_word763_in;
  logic [64:0] zll_main_word764_in;
  logic [63:0] zll_main_word767_in;
  logic [63:0] zll_main_word766_in;
  logic [71:0] zll_pure_dispatch91_in;
  logic [64:0] main_word85_in;
  logic [97:0] zll_main_word854_in;
  logic [64:0] zll_main_word852_in;
  logic [64:0] zll_main_word85_in;
  logic [31:0] zll_main_word856_in;
  logic [64:0] zll_main_word855_in;
  logic [63:0] zll_main_word853_in;
  logic [63:0] zll_main_word851_in;
  logic [71:0] zll_pure_dispatch122_in;
  logic [64:0] main_word91_in;
  logic [97:0] zll_main_word91_in;
  logic [64:0] zll_main_word913_in;
  logic [64:0] zll_main_word912_in;
  logic [31:0] zll_main_word915_in;
  logic [64:0] zll_main_word911_in;
  logic [63:0] zll_main_word914_in;
  logic [63:0] zll_main_word916_in;
  logic [71:0] zll_pure_dispatch13_in;
  logic [64:0] main_word5_in;
  logic [97:0] zll_main_word515_in;
  logic [64:0] zll_main_word527_in;
  logic [64:0] zll_main_word519_in;
  logic [31:0] zll_main_word517_in;
  logic [64:0] zll_main_word528_in;
  logic [63:0] zll_main_word54_in;
  logic [63:0] zll_main_word513_in;
  logic [63:0] zll_main_word430_inR2;
  logic [65:0] zll_main_word430_outR2;
  logic [97:0] zll_main_word5_in;
  logic [97:0] zll_main_word530_in;
  logic [95:0] zll_main_word514_in;
  logic [63:0] test3_in;
  logic [0:0] extresR2;
  logic [71:0] zll_pure_dispatch6_in;
  logic [64:0] main_word75_in;
  logic [97:0] zll_main_word755_in;
  logic [64:0] zll_main_word756_in;
  logic [64:0] zll_main_word754_in;
  logic [31:0] zll_main_word75_in;
  logic [64:0] zll_main_word753_in;
  logic [63:0] zll_main_word752_in;
  logic [63:0] zll_main_word751_in;
  logic [71:0] zll_pure_dispatch66_in;
  logic [64:0] main_word86_in;
  logic [97:0] zll_main_word862_in;
  logic [64:0] zll_main_word861_in;
  logic [64:0] zll_main_word865_in;
  logic [31:0] zll_main_word864_in;
  logic [64:0] zll_main_word86_in;
  logic [63:0] zll_main_word866_in;
  logic [63:0] zll_main_word863_in;
  logic [71:0] zll_pure_dispatch17_in;
  logic [64:0] main_word7_in;
  logic [97:0] zll_main_word7_in;
  logic [64:0] zll_main_word717_in;
  logic [64:0] zll_main_word720_in;
  logic [31:0] zll_main_word715_in;
  logic [64:0] zll_main_word710_in;
  logic [63:0] zll_main_word76_in;
  logic [63:0] zll_main_word714_in;
  logic [71:0] zll_pure_dispatch63_in;
  logic [64:0] main_word3_in;
  logic [97:0] zll_main_word337_in;
  logic [64:0] zll_main_word310_in;
  logic [64:0] zll_main_word314_in;
  logic [65:0] zll_main_word314_out;
  logic [64:0] zll_main_word37_in;
  logic [63:0] zll_main_word313_in;
  logic [63:0] zll_main_word317_in;
  logic [63:0] zll_main_word430_inR3;
  logic [65:0] zll_main_word430_outR3;
  logic [97:0] zll_main_word33_in;
  logic [97:0] zll_main_word329_in;
  logic [95:0] zll_main_word3_in;
  logic [63:0] test1_inR1;
  logic [0:0] extresR3;
  logic [71:0] zll_pure_dispatch112_in;
  logic [64:0] main_word45_in;
  logic [97:0] zll_main_word456_in;
  logic [64:0] zll_main_word45_in;
  logic [64:0] zll_main_word455_in;
  logic [31:0] zll_main_word453_in;
  logic [64:0] zll_main_word451_in;
  logic [63:0] zll_main_word452_in;
  logic [63:0] zll_main_word454_in;
  logic [71:0] zll_pure_dispatch26_in;
  logic [64:0] main_word43_in;
  logic [97:0] zll_main_word433_in;
  logic [64:0] zll_main_word435_in;
  logic [64:0] zll_main_word437_in;
  logic [31:0] zll_main_word432_in;
  logic [64:0] zll_main_word431_in;
  logic [63:0] zll_main_word434_in;
  logic [63:0] zll_main_word436_in;
  logic [71:0] zll_pure_dispatch_in;
  logic [64:0] main_word116_in;
  logic [97:0] zll_main_word1166_in;
  logic [64:0] zll_main_word1167_in;
  logic [64:0] zll_main_word1165_in;
  logic [31:0] zll_main_word1162_in;
  logic [64:0] zll_main_word1161_in;
  logic [63:0] zll_main_word1164_in;
  logic [63:0] zll_main_word1163_in;
  logic [71:0] zll_pure_dispatch118_in;
  logic [64:0] main_word54_in;
  logic [97:0] zll_main_word541_in;
  logic [64:0] zll_main_word547_in;
  logic [64:0] zll_main_word543_in;
  logic [31:0] zll_main_word542_in;
  logic [64:0] zll_main_word545_in;
  logic [63:0] zll_main_word546_in;
  logic [63:0] zll_main_word544_in;
  logic [71:0] zll_pure_dispatch126_in;
  logic [64:0] main_word113_in;
  logic [97:0] zll_main_word1135_in;
  logic [64:0] zll_main_word1134_in;
  logic [64:0] zll_main_word1136_in;
  logic [31:0] zll_main_word1132_in;
  logic [64:0] zll_main_word1131_in;
  logic [63:0] zll_main_word1133_in;
  logic [63:0] zll_main_word113_in;
  logic [71:0] zll_pure_dispatch83_in;
  logic [64:0] main_word47_in;
  logic [97:0] zll_main_word474_in;
  logic [64:0] zll_main_word471_in;
  logic [64:0] zll_main_word473_in;
  logic [31:0] zll_main_word47_in;
  logic [64:0] zll_main_word476_in;
  logic [63:0] zll_main_word472_in;
  logic [63:0] zll_main_word475_in;
  logic [71:0] zll_pure_dispatch102_in;
  logic [64:0] main_word60_in;
  logic [97:0] zll_main_word606_in;
  logic [64:0] zll_main_word60_in;
  logic [64:0] zll_main_word603_in;
  logic [31:0] zll_main_word604_in;
  logic [64:0] zll_main_word605_in;
  logic [63:0] zll_main_word602_in;
  logic [63:0] zll_main_word601_in;
  logic [71:0] zll_pure_dispatch33_in;
  logic [64:0] main_word72_in;
  logic [97:0] zll_main_word725_in;
  logic [64:0] zll_main_word72_in;
  logic [64:0] zll_main_word721_in;
  logic [31:0] zll_main_word723_in;
  logic [64:0] zll_main_word722_in;
  logic [63:0] zll_main_word726_in;
  logic [63:0] zll_main_word724_in;
  logic [71:0] zll_pure_dispatch50_in;
  logic [64:0] main_word79_in;
  logic [97:0] zll_main_word791_in;
  logic [64:0] zll_main_word796_in;
  logic [64:0] zll_main_word79_in;
  logic [31:0] zll_main_word795_in;
  logic [64:0] zll_main_word794_in;
  logic [63:0] zll_main_word793_in;
  logic [63:0] zll_main_word792_in;
  logic [71:0] zll_pure_dispatch56_in;
  logic [64:0] main_word6_in;
  logic [97:0] zll_main_word65_in;
  logic [64:0] zll_main_word629_in;
  logic [64:0] zll_main_word610_in;
  logic [31:0] zll_main_word611_in;
  logic [64:0] zll_main_word617_in;
  logic [63:0] zll_main_word619_in;
  logic [63:0] zll_main_word6_in;
  logic [63:0] zll_main_word430_inR4;
  logic [65:0] zll_main_word430_outR4;
  logic [97:0] zll_main_word626_in;
  logic [97:0] zll_main_word625_in;
  logic [95:0] zll_main_word620_in;
  logic [63:0] test4_in;
  logic [0:0] extresR4;
  logic [71:0] zll_pure_dispatch47_in;
  logic [64:0] main_word74_in;
  logic [97:0] zll_main_word745_in;
  logic [64:0] zll_main_word74_in;
  logic [64:0] zll_main_word744_in;
  logic [31:0] zll_main_word743_in;
  logic [64:0] zll_main_word746_in;
  logic [63:0] zll_main_word741_in;
  logic [63:0] zll_main_word742_in;
  logic [71:0] zll_pure_dispatch53_in;
  logic [64:0] main_word28_in;
  logic [97:0] zll_main_word282_in;
  logic [64:0] zll_main_word283_in;
  logic [64:0] zll_main_word28_in;
  logic [31:0] zll_main_word281_in;
  logic [64:0] zll_main_word286_in;
  logic [63:0] zll_main_word284_in;
  logic [63:0] zll_main_word285_in;
  logic [71:0] zll_pure_dispatch31_in;
  logic [64:0] main_word38_in;
  logic [97:0] zll_main_word385_in;
  logic [64:0] zll_main_word384_in;
  logic [64:0] zll_main_word386_in;
  logic [31:0] zll_main_word383_in;
  logic [64:0] zll_main_word382_in;
  logic [63:0] zll_main_word38_in;
  logic [63:0] zll_main_word381_in;
  logic [71:0] zll_pure_dispatch25_in;
  logic [64:0] main_word15_in;
  logic [97:0] zll_main_word156_in;
  logic [64:0] zll_main_word155_in;
  logic [64:0] zll_main_word151_in;
  logic [31:0] zll_main_word153_in;
  logic [64:0] zll_main_word154_in;
  logic [63:0] zll_main_word152_in;
  logic [63:0] zll_main_word15_in;
  logic [71:0] zll_pure_dispatch115_in;
  logic [64:0] main_word99_in;
  logic [97:0] zll_main_word993_in;
  logic [64:0] zll_main_word996_in;
  logic [64:0] zll_main_word994_in;
  logic [31:0] zll_main_word991_in;
  logic [64:0] zll_main_word995_in;
  logic [63:0] zll_main_word992_in;
  logic [63:0] zll_main_word99_in;
  logic [71:0] zll_pure_dispatch11_in;
  logic [64:0] main_word20_in;
  logic [97:0] zll_main_word204_in;
  logic [64:0] zll_main_word202_in;
  logic [64:0] zll_main_word201_in;
  logic [31:0] zll_main_word205_in;
  logic [64:0] zll_main_word20_in;
  logic [63:0] zll_main_word203_in;
  logic [63:0] zll_main_word206_in;
  logic [71:0] zll_pure_dispatch101_in;
  logic [64:0] main_word9_in;
  logic [97:0] zll_main_word9_in;
  logic [64:0] zll_main_word917_in;
  logic [64:0] zll_main_word910_in;
  logic [31:0] zll_main_word92_in;
  logic [64:0] zll_main_word918_in;
  logic [63:0] zll_main_word919_in;
  logic [63:0] zll_main_word920_in;
  logic [71:0] zll_pure_dispatch18_in;
  logic [64:0] main_word14_in;
  logic [97:0] zll_main_word142_in;
  logic [64:0] zll_main_word148_in;
  logic [64:0] zll_main_word143_in;
  logic [31:0] zll_main_word146_in;
  logic [64:0] zll_main_word141_in;
  logic [63:0] zll_main_word144_in;
  logic [63:0] zll_main_word145_in;
  logic [71:0] zll_pure_dispatch81_in;
  logic [64:0] main_word29_in;
  logic [97:0] zll_main_word295_in;
  logic [64:0] zll_main_word291_in;
  logic [64:0] zll_main_word292_in;
  logic [31:0] zll_main_word29_in;
  logic [64:0] zll_main_word293_in;
  logic [63:0] zll_main_word296_in;
  logic [63:0] zll_main_word294_in;
  logic [71:0] zll_pure_dispatch108_in;
  logic [64:0] main_word95_in;
  logic [97:0] zll_main_word953_in;
  logic [64:0] zll_main_word955_in;
  logic [64:0] zll_main_word954_in;
  logic [31:0] zll_main_word95_in;
  logic [64:0] zll_main_word952_in;
  logic [63:0] zll_main_word956_in;
  logic [63:0] zll_main_word951_in;
  logic [71:0] zll_pure_dispatch46_in;
  logic [64:0] main_word77_in;
  logic [97:0] zll_main_word776_in;
  logic [64:0] zll_main_word77_in;
  logic [64:0] zll_main_word773_in;
  logic [31:0] zll_main_word772_in;
  logic [64:0] zll_main_word774_in;
  logic [63:0] zll_main_word771_in;
  logic [63:0] zll_main_word775_in;
  logic [71:0] zll_pure_dispatch104_in;
  logic [64:0] main_word119_in;
  logic [97:0] zll_main_word1195_in;
  logic [64:0] zll_main_word1196_in;
  logic [64:0] zll_main_word1191_in;
  logic [31:0] zll_main_word119_in;
  logic [64:0] zll_main_word1192_in;
  logic [63:0] zll_main_word1193_in;
  logic [63:0] zll_main_word1194_in;
  logic [71:0] zll_pure_dispatch3_in;
  logic [64:0] main_word63_in;
  logic [97:0] zll_main_word631_in;
  logic [64:0] zll_main_word634_in;
  logic [64:0] zll_main_word633_in;
  logic [31:0] zll_main_word635_in;
  logic [64:0] zll_main_word63_in;
  logic [63:0] zll_main_word636_in;
  logic [63:0] zll_main_word632_in;
  logic [71:0] zll_pure_dispatch38_in;
  logic [64:0] main_word65_in;
  logic [97:0] zll_main_word654_in;
  logic [64:0] zll_main_word653_in;
  logic [64:0] zll_main_word656_in;
  logic [31:0] zll_main_word657_in;
  logic [64:0] zll_main_word655_in;
  logic [63:0] zll_main_word651_in;
  logic [63:0] zll_main_word652_in;
  logic [71:0] zll_pure_dispatch78_in;
  logic [64:0] main_word78_in;
  logic [97:0] zll_main_word78_in;
  logic [64:0] zll_main_word785_in;
  logic [64:0] zll_main_word786_in;
  logic [31:0] zll_main_word783_in;
  logic [64:0] zll_main_word782_in;
  logic [63:0] zll_main_word784_in;
  logic [63:0] zll_main_word781_in;
  logic [71:0] zll_pure_dispatch89_in;
  logic [64:0] main_word57_in;
  logic [97:0] zll_main_word574_in;
  logic [64:0] zll_main_word571_in;
  logic [64:0] zll_main_word573_in;
  logic [31:0] zll_main_word575_in;
  logic [64:0] zll_main_word57_in;
  logic [63:0] zll_main_word572_in;
  logic [63:0] zll_main_word576_in;
  logic [71:0] zll_pure_dispatch14_in;
  logic [64:0] main_word121_in;
  logic [97:0] zll_main_word12111_in;
  logic [64:0] zll_main_word1214_in;
  logic [64:0] zll_main_word1212_in;
  logic [31:0] zll_main_word12110_in;
  logic [64:0] zll_main_word1217_in;
  logic [63:0] zll_main_word1216_in;
  logic [63:0] zll_main_word1218_in;
  logic [71:0] zll_pure_dispatch106_in;
  logic [64:0] main_word40_in;
  logic [97:0] zll_main_word40_in;
  logic [64:0] zll_main_word403_in;
  logic [64:0] zll_main_word402_in;
  logic [31:0] zll_main_word404_in;
  logic [64:0] zll_main_word401_in;
  logic [63:0] zll_main_word406_in;
  logic [63:0] zll_main_word405_in;
  logic [71:0] zll_pure_dispatch70_in;
  logic [64:0] main_word67_in;
  logic [97:0] zll_main_word671_in;
  logic [64:0] zll_main_word673_in;
  logic [64:0] zll_main_word676_in;
  logic [31:0] zll_main_word67_in;
  logic [64:0] zll_main_word674_in;
  logic [63:0] zll_main_word675_in;
  logic [63:0] zll_main_word672_in;
  logic [71:0] zll_pure_dispatch39_in;
  logic [64:0] main_word33_in;
  logic [97:0] zll_main_word335_in;
  logic [64:0] zll_main_word338_in;
  logic [64:0] zll_main_word332_in;
  logic [31:0] zll_main_word336_in;
  logic [64:0] zll_main_word334_in;
  logic [63:0] zll_main_word333_in;
  logic [63:0] zll_main_word331_in;
  logic [71:0] zll_pure_dispatch84_in;
  logic [64:0] main_word22_in;
  logic [97:0] zll_main_word228_in;
  logic [64:0] zll_main_word223_in;
  logic [64:0] zll_main_word222_in;
  logic [31:0] zll_main_word229_in;
  logic [64:0] zll_main_word22_in;
  logic [63:0] zll_main_word224_in;
  logic [63:0] zll_main_word221_in;
  logic [71:0] zll_pure_dispatch60_in;
  logic [64:0] main_word93_in;
  logic [97:0] zll_main_word932_in;
  logic [64:0] zll_main_word933_in;
  logic [64:0] zll_main_word934_in;
  logic [31:0] zll_main_word93_in;
  logic [64:0] zll_main_word935_in;
  logic [63:0] zll_main_word931_in;
  logic [63:0] zll_main_word936_in;
  logic [71:0] zll_pure_dispatch105_in;
  logic [64:0] main_word36_in;
  logic [97:0] zll_main_word365_in;
  logic [64:0] zll_main_word362_in;
  logic [64:0] zll_main_word361_in;
  logic [31:0] zll_main_word366_in;
  logic [64:0] zll_main_word36_in;
  logic [63:0] zll_main_word363_in;
  logic [63:0] zll_main_word364_in;
  logic [71:0] zll_pure_dispatch107_in;
  logic [64:0] main_word110_in;
  logic [97:0] zll_main_word1105_in;
  logic [64:0] zll_main_word1103_in;
  logic [64:0] zll_main_word1102_in;
  logic [31:0] zll_main_word1104_in;
  logic [64:0] zll_main_word110_in;
  logic [63:0] zll_main_word1106_in;
  logic [63:0] zll_main_word1101_in;
  logic [71:0] zll_pure_dispatch109_in;
  logic [64:0] main_word84_in;
  logic [97:0] zll_main_word841_in;
  logic [64:0] zll_main_word844_in;
  logic [64:0] zll_main_word846_in;
  logic [31:0] zll_main_word843_in;
  logic [64:0] zll_main_word845_in;
  logic [63:0] zll_main_word842_in;
  logic [63:0] zll_main_word84_in;
  logic [71:0] zll_pure_dispatch4_in;
  logic [64:0] main_word97_in;
  logic [97:0] zll_main_word976_in;
  logic [64:0] zll_main_word973_in;
  logic [64:0] zll_main_word974_in;
  logic [31:0] zll_main_word97_in;
  logic [64:0] zll_main_word972_in;
  logic [63:0] zll_main_word971_in;
  logic [63:0] zll_main_word975_in;
  logic [71:0] zll_pure_dispatch61_in;
  logic [64:0] main_word11_in;
  logic [97:0] zll_main_word1114_in;
  logic [64:0] zll_main_word1116_in;
  logic [64:0] zll_main_word1117_in;
  logic [31:0] zll_main_word1110_in;
  logic [64:0] zll_main_word1120_in;
  logic [63:0] zll_main_word11_in;
  logic [63:0] zll_main_word116_in;
  logic [71:0] zll_pure_dispatch16_in;
  logic [64:0] main_word88_in;
  logic [97:0] zll_main_word885_in;
  logic [64:0] zll_main_word886_in;
  logic [64:0] zll_main_word884_in;
  logic [31:0] zll_main_word881_in;
  logic [64:0] zll_main_word88_in;
  logic [63:0] zll_main_word883_in;
  logic [63:0] zll_main_word882_in;
  logic [71:0] zll_pure_dispatch51_in;
  logic [64:0] main_word46_in;
  logic [97:0] zll_main_word46_in;
  logic [64:0] zll_main_word464_in;
  logic [64:0] zll_main_word461_in;
  logic [31:0] zll_main_word466_in;
  logic [64:0] zll_main_word462_in;
  logic [63:0] zll_main_word463_in;
  logic [63:0] zll_main_word465_in;
  logic [71:0] zll_pure_dispatch24_in;
  logic [64:0] main_word105_in;
  logic [97:0] zll_main_word1054_in;
  logic [64:0] zll_main_word1052_in;
  logic [64:0] zll_main_word1053_in;
  logic [31:0] zll_main_word1051_in;
  logic [64:0] zll_main_word1055_in;
  logic [63:0] zll_main_word105_in;
  logic [63:0] zll_main_word1056_in;
  logic [71:0] zll_pure_dispatch119_in;
  logic [64:0] main_word01_in;
  logic [97:0] zll_main_word012_in;
  logic [64:0] zll_main_word011_in;
  logic [64:0] zll_main_word010_in;
  logic [31:0] zll_main_word08_in;
  logic [64:0] zll_main_word01_in;
  logic [63:0] zll_main_word07_in;
  logic [63:0] zll_main_word04_in;
  logic [31:0] zll_main_word06_in;
  logic [65:0] zll_main_word06_out;
  logic [65:0] zll_main_word05_in;
  logic [65:0] zll_main_word09_inR1;
  logic [65:0] zll_main_word09_outR1;
  logic [71:0] zll_pure_dispatch65_in;
  logic [64:0] main_word62_in;
  logic [97:0] zll_main_word62_in;
  logic [64:0] zll_main_word627_in;
  logic [64:0] zll_main_word621_in;
  logic [31:0] zll_main_word628_in;
  logic [64:0] zll_main_word624_in;
  logic [63:0] zll_main_word623_in;
  logic [63:0] zll_main_word622_in;
  logic [71:0] zll_pure_dispatch55_in;
  logic [64:0] main_word2_in;
  logic [97:0] zll_main_word226_in;
  logic [64:0] zll_main_word225_in;
  logic [64:0] zll_main_word227_in;
  logic [31:0] zll_main_word230_in;
  logic [64:0] zll_main_word220_in;
  logic [63:0] zll_main_word214_in;
  logic [63:0] zll_main_word21_in;
  logic [31:0] zll_main_word06_inR1;
  logic [65:0] zll_main_word06_outR1;
  logic [65:0] zll_main_word211_in;
  logic [65:0] zll_main_word314_inR1;
  logic [65:0] zll_main_word314_outR1;
  logic [71:0] zll_pure_dispatch125_in;
  logic [64:0] main_word30_in;
  logic [97:0] zll_main_word301_in;
  logic [64:0] zll_main_word302_in;
  logic [64:0] zll_main_word304_in;
  logic [31:0] zll_main_word30_in;
  logic [64:0] zll_main_word305_in;
  logic [63:0] zll_main_word303_in;
  logic [63:0] zll_main_word306_in;
  logic [71:0] zll_pure_dispatch98_in;
  logic [64:0] main_word90_in;
  logic [97:0] zll_main_word90_in;
  logic [64:0] zll_main_word902_in;
  logic [64:0] zll_main_word905_in;
  logic [31:0] zll_main_word901_in;
  logic [64:0] zll_main_word906_in;
  logic [63:0] zll_main_word904_in;
  logic [63:0] zll_main_word903_in;
  logic [71:0] zll_pure_dispatch29_in;
  logic [64:0] main_word109_in;
  logic [97:0] zll_main_word109_in;
  logic [64:0] zll_main_word1093_in;
  logic [64:0] zll_main_word1091_in;
  logic [31:0] zll_main_word1095_in;
  logic [64:0] zll_main_word1094_in;
  logic [63:0] zll_main_word1096_in;
  logic [63:0] zll_main_word1092_in;
  logic [71:0] zll_pure_dispatch100_in;
  logic [64:0] main_word34_in;
  logic [97:0] zll_main_word344_in;
  logic [64:0] zll_main_word342_in;
  logic [64:0] zll_main_word343_in;
  logic [31:0] zll_main_word341_in;
  logic [64:0] zll_main_word346_in;
  logic [63:0] zll_main_word345_in;
  logic [63:0] zll_main_word34_in;
  logic [71:0] zll_pure_dispatch121_in;
  logic [64:0] main_word108_in;
  logic [97:0] zll_main_word1082_in;
  logic [64:0] zll_main_word1085_in;
  logic [64:0] zll_main_word1086_in;
  logic [31:0] zll_main_word1087_in;
  logic [64:0] zll_main_word1083_in;
  logic [63:0] zll_main_word1081_in;
  logic [63:0] zll_main_word1084_in;
  logic [71:0] zll_pure_dispatch40_in;
  logic [64:0] main_word44_in;
  logic [97:0] zll_main_word44_in;
  logic [64:0] zll_main_word446_in;
  logic [64:0] zll_main_word441_in;
  logic [31:0] zll_main_word444_in;
  logic [64:0] zll_main_word445_in;
  logic [63:0] zll_main_word442_in;
  logic [63:0] zll_main_word443_in;
  logic [71:0] zll_pure_dispatch30_in;
  logic [64:0] main_word64_in;
  logic [97:0] zll_main_word641_in;
  logic [64:0] zll_main_word643_in;
  logic [64:0] zll_main_word642_in;
  logic [31:0] zll_main_word645_in;
  logic [64:0] zll_main_word646_in;
  logic [63:0] zll_main_word644_in;
  logic [63:0] zll_main_word647_in;
  logic [71:0] zll_pure_dispatch120_in;
  logic [64:0] main_word49_in;
  logic [97:0] zll_main_word496_in;
  logic [64:0] zll_main_word491_in;
  logic [64:0] zll_main_word495_in;
  logic [31:0] zll_main_word494_in;
  logic [64:0] zll_main_word49_in;
  logic [63:0] zll_main_word492_in;
  logic [63:0] zll_main_word493_in;
  logic [71:0] zll_pure_dispatch73_in;
  logic [64:0] main_word73_in;
  logic [97:0] zll_main_word73_in;
  logic [64:0] zll_main_word734_in;
  logic [64:0] zll_main_word733_in;
  logic [31:0] zll_main_word736_in;
  logic [64:0] zll_main_word735_in;
  logic [63:0] zll_main_word731_in;
  logic [63:0] zll_main_word732_in;
  logic [71:0] zll_pure_dispatch23_in;
  logic [64:0] main_word114_in;
  logic [97:0] zll_main_word1141_in;
  logic [64:0] zll_main_word1144_in;
  logic [64:0] zll_main_word1145_in;
  logic [31:0] zll_main_word1146_in;
  logic [64:0] zll_main_word1143_in;
  logic [63:0] zll_main_word114_in;
  logic [63:0] zll_main_word1142_in;
  logic [71:0] zll_pure_dispatch43_in;
  logic [64:0] main_word124_in;
  logic [97:0] zll_main_word1243_in;
  logic [64:0] zll_main_word1247_in;
  logic [64:0] zll_main_word1245_in;
  logic [31:0] zll_main_word1246_in;
  logic [64:0] zll_main_word1244_in;
  logic [63:0] zll_main_word1241_in;
  logic [63:0] zll_main_word1242_in;
  logic [71:0] zll_pure_dispatch95_in;
  logic [64:0] main_word48_in;
  logic [97:0] zll_main_word485_in;
  logic [64:0] zll_main_word483_in;
  logic [64:0] zll_main_word486_in;
  logic [31:0] zll_main_word481_in;
  logic [64:0] zll_main_word48_in;
  logic [63:0] zll_main_word482_in;
  logic [63:0] zll_main_word484_in;
  logic [71:0] zll_pure_dispatch75_in;
  logic [64:0] main_word117_in;
  logic [97:0] zll_main_word1172_in;
  logic [64:0] zll_main_word1175_in;
  logic [64:0] zll_main_word1176_in;
  logic [31:0] zll_main_word1173_in;
  logic [64:0] zll_main_word117_in;
  logic [63:0] zll_main_word1171_in;
  logic [63:0] zll_main_word1174_in;
  logic [71:0] zll_pure_dispatch52_in;
  logic [64:0] main_word92_in;
  logic [97:0] zll_main_word925_in;
  logic [64:0] zll_main_word927_in;
  logic [64:0] zll_main_word924_in;
  logic [31:0] zll_main_word922_in;
  logic [64:0] zll_main_word921_in;
  logic [63:0] zll_main_word926_in;
  logic [63:0] zll_main_word923_in;
  logic [71:0] zll_pure_dispatch28_in;
  logic [64:0] main_word120_in;
  logic [97:0] zll_main_word1202_in;
  logic [64:0] zll_main_word1201_in;
  logic [64:0] zll_main_word1204_in;
  logic [31:0] zll_main_word120_in;
  logic [64:0] zll_main_word1205_in;
  logic [63:0] zll_main_word1203_in;
  logic [63:0] zll_main_word1206_in;
  logic [71:0] zll_pure_dispatch59_in;
  logic [64:0] main_word104_in;
  logic [97:0] zll_main_word104_in;
  logic [64:0] zll_main_word1042_in;
  logic [64:0] zll_main_word1044_in;
  logic [31:0] zll_main_word1043_in;
  logic [64:0] zll_main_word1045_in;
  logic [63:0] zll_main_word1046_in;
  logic [63:0] zll_main_word1041_in;
  logic [71:0] zll_pure_dispatch113_in;
  logic [64:0] main_word8_in;
  logic [97:0] zll_main_word82_in;
  logic [64:0] zll_main_word81_in;
  logic [64:0] zll_main_word820_in;
  logic [31:0] zll_main_word815_in;
  logic [64:0] zll_main_word810_in;
  logic [63:0] zll_main_word819_in;
  logic [63:0] zll_main_word8_in;
  logic [71:0] zll_pure_dispatch67_in;
  logic [64:0] main_word17_in;
  logic [97:0] zll_main_word174_in;
  logic [64:0] zll_main_word175_in;
  logic [64:0] zll_main_word176_in;
  logic [31:0] zll_main_word173_in;
  logic [64:0] zll_main_word17_in;
  logic [63:0] zll_main_word172_in;
  logic [63:0] zll_main_word171_in;
  logic [71:0] zll_pure_dispatch36_in;
  logic [64:0] main_word50_in;
  logic [97:0] zll_main_word506_in;
  logic [64:0] zll_main_word502_in;
  logic [64:0] zll_main_word505_in;
  logic [31:0] zll_main_word504_in;
  logic [64:0] zll_main_word501_in;
  logic [63:0] zll_main_word503_in;
  logic [63:0] zll_main_word50_in;
  logic [71:0] zll_pure_dispatch34_in;
  logic [64:0] main_word56_in;
  logic [97:0] zll_main_word56_in;
  logic [64:0] zll_main_word561_in;
  logic [64:0] zll_main_word562_in;
  logic [31:0] zll_main_word564_in;
  logic [64:0] zll_main_word566_in;
  logic [63:0] zll_main_word565_in;
  logic [63:0] zll_main_word563_in;
  logic [71:0] zll_pure_dispatch2_in;
  logic [64:0] main_word70_in;
  logic [97:0] zll_main_word706_in;
  logic [64:0] zll_main_word701_in;
  logic [64:0] zll_main_word704_in;
  logic [31:0] zll_main_word70_in;
  logic [64:0] zll_main_word703_in;
  logic [63:0] zll_main_word702_in;
  logic [63:0] zll_main_word705_in;
  logic [71:0] zll_pure_dispatch54_in;
  logic [64:0] main_word106_in;
  logic [97:0] zll_main_word1061_in;
  logic [64:0] zll_main_word1062_in;
  logic [64:0] zll_main_word1066_in;
  logic [31:0] zll_main_word1064_in;
  logic [64:0] zll_main_word1065_in;
  logic [63:0] zll_main_word106_in;
  logic [63:0] zll_main_word1063_in;
  logic [71:0] zll_pure_dispatch1_in;
  logic [64:0] main_word66_in;
  logic [97:0] zll_main_word667_in;
  logic [64:0] zll_main_word661_in;
  logic [64:0] zll_main_word663_in;
  logic [31:0] zll_main_word665_in;
  logic [64:0] zll_main_word664_in;
  logic [63:0] zll_main_word662_in;
  logic [63:0] zll_main_word666_in;
  logic [71:0] zll_pure_dispatch35_in;
  logic [64:0] main_word23_in;
  logic [97:0] zll_main_word235_in;
  logic [64:0] zll_main_word234_in;
  logic [64:0] zll_main_word236_in;
  logic [31:0] zll_main_word232_in;
  logic [64:0] zll_main_word233_in;
  logic [63:0] zll_main_word231_in;
  logic [63:0] zll_main_word23_in;
  logic [0:0] __continue;
  logic [23:0] __padding;
  logic [6:0] __resumption_tag;
  logic [31:0] __st0;
  logic [6:0] __resumption_tag_next;
  logic [31:0] __st0_next;
  assign zll_pure_dispatch22_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word102_in = {zll_pure_dispatch22_in[71:39], zll_pure_dispatch22_in[31:0]};
  assign zll_main_word1026_in = {main_word102_in[64:32], main_word102_in[64:32], main_word102_in[31:0]};
  assign zll_main_word1023_in = {zll_main_word1026_in[97:65], zll_main_word1026_in[31:0]};
  assign zll_main_word1024_in = {zll_main_word1023_in[31:0], zll_main_word1023_in[64:32]};
  assign zll_main_word1021_in = zll_main_word1024_in[64:33];
  assign zll_main_word102_in = {zll_main_word1026_in[31:0], zll_main_word1026_in[64:32]};
  assign zll_main_word1022_in = {zll_main_word102_in[64:33], zll_main_word102_in[31:0]};
  assign zll_main_word1025_in = {zll_main_word1022_in[31:0], zll_main_word1022_in[63:32]};
  assign zll_pure_dispatch74_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word24_in = {zll_pure_dispatch74_in[71:39], zll_pure_dispatch74_in[31:0]};
  assign zll_main_word246_in = {main_word24_in[64:32], main_word24_in[64:32], main_word24_in[31:0]};
  assign zll_main_word24_in = {zll_main_word246_in[97:65], zll_main_word246_in[31:0]};
  assign zll_main_word245_in = {zll_main_word24_in[31:0], zll_main_word24_in[64:32]};
  assign zll_main_word244_in = zll_main_word245_in[64:33];
  assign zll_main_word241_in = {zll_main_word246_in[31:0], zll_main_word246_in[64:32]};
  assign zll_main_word242_in = {zll_main_word241_in[64:33], zll_main_word241_in[31:0]};
  assign zll_main_word243_in = {zll_main_word242_in[31:0], zll_main_word242_in[63:32]};
  assign zll_pure_dispatch20_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word111_in = {zll_pure_dispatch20_in[71:39], zll_pure_dispatch20_in[31:0]};
  assign zll_main_word1115_in = {main_word111_in[64:32], main_word111_in[64:32], main_word111_in[31:0]};
  assign zll_main_word1113_in = {zll_main_word1115_in[97:65], zll_main_word1115_in[31:0]};
  assign zll_main_word111_in = {zll_main_word1113_in[31:0], zll_main_word1113_in[64:32]};
  assign zll_main_word1119_in = zll_main_word111_in[64:33];
  assign zll_main_word1118_in = {zll_main_word1115_in[31:0], zll_main_word1115_in[64:32]};
  assign zll_main_word1112_in = {zll_main_word1118_in[64:33], zll_main_word1118_in[31:0]};
  assign zll_main_word1111_in = {zll_main_word1112_in[31:0], zll_main_word1112_in[63:32]};
  assign zll_pure_dispatch94_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word10_in = {zll_pure_dispatch94_in[71:39], zll_pure_dispatch94_in[31:0]};
  assign zll_main_word1018_in = {main_word10_in[64:32], main_word10_in[64:32], main_word10_in[31:0]};
  assign zll_main_word108_in = {zll_main_word1018_in[97:65], zll_main_word1018_in[31:0]};
  assign zll_main_word1010_in = {zll_main_word108_in[31:0], zll_main_word108_in[64:32]};
  assign zll_main_word10_in = zll_main_word1010_in[64:33];
  assign zll_main_word1015_in = {zll_main_word1018_in[31:0], zll_main_word1018_in[64:32]};
  assign zll_main_word101_in = {zll_main_word1015_in[64:33], zll_main_word1015_in[31:0]};
  assign zll_main_word1017_in = {zll_main_word101_in[31:0], zll_main_word101_in[63:32]};
  assign zll_pure_dispatch5_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word51_in = {zll_pure_dispatch5_in[71:39], zll_pure_dispatch5_in[31:0]};
  assign zll_main_word511_in = {main_word51_in[64:32], main_word51_in[64:32], main_word51_in[31:0]};
  assign zll_main_word518_in = {zll_main_word511_in[97:65], zll_main_word511_in[31:0]};
  assign zll_main_word516_in = {zll_main_word518_in[31:0], zll_main_word518_in[64:32]};
  assign zll_main_word5111_in = zll_main_word516_in[64:33];
  assign zll_main_word5110_in = {zll_main_word511_in[31:0], zll_main_word511_in[64:32]};
  assign zll_main_word512_in = {zll_main_word5110_in[64:33], zll_main_word5110_in[31:0]};
  assign zll_main_word51_in = {zll_main_word512_in[31:0], zll_main_word512_in[63:32]};
  assign zll_pure_dispatch45_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word4_in = {zll_pure_dispatch45_in[71:39], zll_pure_dispatch45_in[31:0]};
  assign zll_main_word420_in = {main_word4_in[64:32], main_word4_in[64:32], main_word4_in[31:0]};
  assign zll_main_word41_in = {zll_main_word420_in[97:65], zll_main_word420_in[31:0]};
  assign zll_main_word425_in = {zll_main_word41_in[31:0], zll_main_word41_in[64:32]};
  assign zll_main_word4_in = zll_main_word425_in[64:33];
  assign zll_main_word423_in = {zll_main_word420_in[31:0], zll_main_word420_in[64:32]};
  assign zll_main_word410_in = {zll_main_word423_in[64:33], zll_main_word423_in[31:0]};
  assign zll_main_word417_in = {zll_main_word410_in[31:0], zll_main_word410_in[63:32]};
  assign zll_main_word430_in = {zll_main_word417_in[31:0], zll_main_word417_in[31:0]};
  ZLL_Main_word430  inst (zll_main_word430_in[63:0], zll_main_word430_out);
  assign zll_main_word43_in = {zll_main_word417_in[63:32], zll_main_word430_out};
  assign zll_main_word428_in = {zll_main_word43_in[97:66], zll_main_word43_in[65:0]};
  assign zll_main_word418_in = {zll_main_word428_in[97:66], zll_main_word428_in[63:32], zll_main_word428_in[31:0]};
  assign test2_in = {zll_main_word418_in[95:64], zll_main_word418_in[63:32]};
  test2  instR1 (test2_in[63:32], test2_in[31:0], extres[0]);
  assign zll_pure_dispatch68_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word71_in = {zll_pure_dispatch68_in[71:39], zll_pure_dispatch68_in[31:0]};
  assign zll_main_word713_in = {main_word71_in[64:32], main_word71_in[64:32], main_word71_in[31:0]};
  assign zll_main_word716_in = {zll_main_word713_in[97:65], zll_main_word713_in[31:0]};
  assign zll_main_word712_in = {zll_main_word716_in[31:0], zll_main_word716_in[64:32]};
  assign zll_main_word71_in = zll_main_word712_in[64:33];
  assign zll_main_word718_in = {zll_main_word713_in[31:0], zll_main_word713_in[64:32]};
  assign zll_main_word711_in = {zll_main_word718_in[64:33], zll_main_word718_in[31:0]};
  assign zll_main_word719_in = {zll_main_word711_in[31:0], zll_main_word711_in[63:32]};
  assign zll_pure_dispatch123_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word103_in = {zll_pure_dispatch123_in[71:39], zll_pure_dispatch123_in[31:0]};
  assign zll_main_word1036_in = {main_word103_in[64:32], main_word103_in[64:32], main_word103_in[31:0]};
  assign zll_main_word103_in = {zll_main_word1036_in[97:65], zll_main_word1036_in[31:0]};
  assign zll_main_word1031_in = {zll_main_word103_in[31:0], zll_main_word103_in[64:32]};
  assign zll_main_word1034_in = zll_main_word1031_in[64:33];
  assign zll_main_word1035_in = {zll_main_word1036_in[31:0], zll_main_word1036_in[64:32]};
  assign zll_main_word1033_in = {zll_main_word1035_in[64:33], zll_main_word1035_in[31:0]};
  assign zll_main_word1032_in = {zll_main_word1033_in[31:0], zll_main_word1033_in[63:32]};
  assign zll_pure_dispatch9_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word122_in = {zll_pure_dispatch9_in[71:39], zll_pure_dispatch9_in[31:0]};
  assign zll_main_word1222_in = {main_word122_in[64:32], main_word122_in[64:32], main_word122_in[31:0]};
  assign zll_main_word1226_in = {zll_main_word1222_in[97:65], zll_main_word1222_in[31:0]};
  assign zll_main_word1225_in = {zll_main_word1226_in[31:0], zll_main_word1226_in[64:32]};
  assign zll_main_word1223_in = zll_main_word1225_in[64:33];
  assign zll_main_word1224_in = {zll_main_word1222_in[31:0], zll_main_word1222_in[64:32]};
  assign zll_main_word1221_in = {zll_main_word1224_in[64:33], zll_main_word1224_in[31:0]};
  assign zll_main_word122_in = {zll_main_word1221_in[31:0], zll_main_word1221_in[63:32]};
  assign zll_pure_dispatch12_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word126_in = {zll_pure_dispatch12_in[71:39], zll_pure_dispatch12_in[31:0]};
  assign zll_main_word1265_in = {main_word126_in[64:32], main_word126_in[64:32], main_word126_in[31:0]};
  assign zll_main_word126_in = {zll_main_word1265_in[97:65], zll_main_word1265_in[31:0]};
  assign zll_main_word1262_in = {zll_main_word126_in[31:0], zll_main_word126_in[64:32]};
  assign zll_main_word1264_in = zll_main_word1262_in[64:33];
  assign zll_main_word1263_in = {zll_main_word1265_in[31:0], zll_main_word1265_in[64:32]};
  assign zll_main_word1261_in = {zll_main_word1263_in[64:33], zll_main_word1263_in[31:0]};
  assign zll_main_word1266_in = {zll_main_word1261_in[31:0], zll_main_word1261_in[63:32]};
  assign zll_pure_dispatch124_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word81_in = {zll_pure_dispatch124_in[71:39], zll_pure_dispatch124_in[31:0]};
  assign zll_main_word813_in = {main_word81_in[64:32], main_word81_in[64:32], main_word81_in[31:0]};
  assign zll_main_word818_in = {zll_main_word813_in[97:65], zll_main_word813_in[31:0]};
  assign zll_main_word812_in = {zll_main_word818_in[31:0], zll_main_word818_in[64:32]};
  assign zll_main_word816_in = zll_main_word812_in[64:33];
  assign zll_main_word811_in = {zll_main_word813_in[31:0], zll_main_word813_in[64:32]};
  assign zll_main_word814_in = {zll_main_word811_in[64:33], zll_main_word811_in[31:0]};
  assign zll_main_word817_in = {zll_main_word814_in[31:0], zll_main_word814_in[63:32]};
  assign zll_pure_dispatch85_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word107_in = {zll_pure_dispatch85_in[71:39], zll_pure_dispatch85_in[31:0]};
  assign zll_main_word1073_in = {main_word107_in[64:32], main_word107_in[64:32], main_word107_in[31:0]};
  assign zll_main_word107_in = {zll_main_word1073_in[97:65], zll_main_word1073_in[31:0]};
  assign zll_main_word1075_in = {zll_main_word107_in[31:0], zll_main_word107_in[64:32]};
  assign zll_main_word1071_in = zll_main_word1075_in[64:33];
  assign zll_main_word1076_in = {zll_main_word1073_in[31:0], zll_main_word1073_in[64:32]};
  assign zll_main_word1072_in = {zll_main_word1076_in[64:33], zll_main_word1076_in[31:0]};
  assign zll_main_word1074_in = {zll_main_word1072_in[31:0], zll_main_word1072_in[63:32]};
  assign zll_pure_dispatch49_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word118_in = {zll_pure_dispatch49_in[71:39], zll_pure_dispatch49_in[31:0]};
  assign zll_main_word1184_in = {main_word118_in[64:32], main_word118_in[64:32], main_word118_in[31:0]};
  assign zll_main_word1182_in = {zll_main_word1184_in[97:65], zll_main_word1184_in[31:0]};
  assign zll_main_word1187_in = {zll_main_word1182_in[31:0], zll_main_word1182_in[64:32]};
  assign zll_main_word1183_in = zll_main_word1187_in[64:33];
  assign zll_main_word1181_in = {zll_main_word1184_in[31:0], zll_main_word1184_in[64:32]};
  assign zll_main_word1185_in = {zll_main_word1181_in[64:33], zll_main_word1181_in[31:0]};
  assign zll_main_word1186_in = {zll_main_word1185_in[31:0], zll_main_word1185_in[63:32]};
  assign zll_pure_dispatch76_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word61_in = {zll_pure_dispatch76_in[71:39], zll_pure_dispatch76_in[31:0]};
  assign zll_main_word616_in = {main_word61_in[64:32], main_word61_in[64:32], main_word61_in[31:0]};
  assign zll_main_word6110_in = {zll_main_word616_in[97:65], zll_main_word616_in[31:0]};
  assign zll_main_word612_in = {zll_main_word6110_in[31:0], zll_main_word6110_in[64:32]};
  assign zll_main_word61_in = zll_main_word612_in[64:33];
  assign zll_main_word6112_in = {zll_main_word616_in[31:0], zll_main_word616_in[64:32]};
  assign zll_main_word618_in = {zll_main_word6112_in[64:33], zll_main_word6112_in[31:0]};
  assign zll_main_word6111_in = {zll_main_word618_in[31:0], zll_main_word618_in[63:32]};
  assign zll_pure_dispatch114_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word98_in = {zll_pure_dispatch114_in[71:39], zll_pure_dispatch114_in[31:0]};
  assign zll_main_word985_in = {main_word98_in[64:32], main_word98_in[64:32], main_word98_in[31:0]};
  assign zll_main_word983_in = {zll_main_word985_in[97:65], zll_main_word985_in[31:0]};
  assign zll_main_word986_in = {zll_main_word983_in[31:0], zll_main_word983_in[64:32]};
  assign zll_main_word98_in = zll_main_word986_in[64:33];
  assign zll_main_word982_in = {zll_main_word985_in[31:0], zll_main_word985_in[64:32]};
  assign zll_main_word981_in = {zll_main_word982_in[64:33], zll_main_word982_in[31:0]};
  assign zll_main_word984_in = {zll_main_word981_in[31:0], zll_main_word981_in[63:32]};
  assign zll_pure_dispatch10_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word18_in = {zll_pure_dispatch10_in[71:39], zll_pure_dispatch10_in[31:0]};
  assign zll_main_word183_in = {main_word18_in[64:32], main_word18_in[64:32], main_word18_in[31:0]};
  assign zll_main_word185_in = {zll_main_word183_in[97:65], zll_main_word183_in[31:0]};
  assign zll_main_word182_in = {zll_main_word185_in[31:0], zll_main_word185_in[64:32]};
  assign zll_main_word18_in = zll_main_word182_in[64:33];
  assign zll_main_word186_in = {zll_main_word183_in[31:0], zll_main_word183_in[64:32]};
  assign zll_main_word184_in = {zll_main_word186_in[64:33], zll_main_word186_in[31:0]};
  assign zll_main_word181_in = {zll_main_word184_in[31:0], zll_main_word184_in[63:32]};
  assign zll_pure_dispatch42_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word100_in = {zll_pure_dispatch42_in[71:39], zll_pure_dispatch42_in[31:0]};
  assign zll_main_word1005_in = {main_word100_in[64:32], main_word100_in[64:32], main_word100_in[31:0]};
  assign zll_main_word1004_in = {zll_main_word1005_in[97:65], zll_main_word1005_in[31:0]};
  assign zll_main_word100_in = {zll_main_word1004_in[31:0], zll_main_word1004_in[64:32]};
  assign zll_main_word1006_in = zll_main_word100_in[64:33];
  assign zll_main_word1003_in = {zll_main_word1005_in[31:0], zll_main_word1005_in[64:32]};
  assign zll_main_word1002_in = {zll_main_word1003_in[64:33], zll_main_word1003_in[31:0]};
  assign zll_main_word1001_in = {zll_main_word1002_in[31:0], zll_main_word1002_in[63:32]};
  assign zll_pure_dispatch37_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word125_in = {zll_pure_dispatch37_in[71:39], zll_pure_dispatch37_in[31:0]};
  assign zll_main_word1254_in = {main_word125_in[64:32], main_word125_in[64:32], main_word125_in[31:0]};
  assign zll_main_word1255_in = {zll_main_word1254_in[97:65], zll_main_word1254_in[31:0]};
  assign zll_main_word1252_in = {zll_main_word1255_in[31:0], zll_main_word1255_in[64:32]};
  assign zll_main_word1251_in = zll_main_word1252_in[64:33];
  assign zll_main_word1256_in = {zll_main_word1254_in[31:0], zll_main_word1254_in[64:32]};
  assign zll_main_word125_in = {zll_main_word1256_in[64:33], zll_main_word1256_in[31:0]};
  assign zll_main_word1253_in = {zll_main_word125_in[31:0], zll_main_word125_in[63:32]};
  assign zll_pure_dispatch96_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word59_in = {zll_pure_dispatch96_in[71:39], zll_pure_dispatch96_in[31:0]};
  assign zll_main_word592_in = {main_word59_in[64:32], main_word59_in[64:32], main_word59_in[31:0]};
  assign zll_main_word596_in = {zll_main_word592_in[97:65], zll_main_word592_in[31:0]};
  assign zll_main_word595_in = {zll_main_word596_in[31:0], zll_main_word596_in[64:32]};
  assign zll_main_word593_in = zll_main_word595_in[64:33];
  assign zll_main_word594_in = {zll_main_word592_in[31:0], zll_main_word592_in[64:32]};
  assign zll_main_word597_in = {zll_main_word594_in[64:33], zll_main_word594_in[31:0]};
  assign zll_main_word591_in = {zll_main_word597_in[31:0], zll_main_word597_in[63:32]};
  assign zll_pure_dispatch99_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word32_in = {zll_pure_dispatch99_in[71:39], zll_pure_dispatch99_in[31:0]};
  assign zll_main_word327_in = {main_word32_in[64:32], main_word32_in[64:32], main_word32_in[31:0]};
  assign zll_main_word324_in = {zll_main_word327_in[97:65], zll_main_word327_in[31:0]};
  assign zll_main_word32_in = {zll_main_word324_in[31:0], zll_main_word324_in[64:32]};
  assign zll_main_word322_in = zll_main_word32_in[64:33];
  assign zll_main_word323_in = {zll_main_word327_in[31:0], zll_main_word327_in[64:32]};
  assign zll_main_word321_in = {zll_main_word323_in[64:33], zll_main_word323_in[31:0]};
  assign zll_main_word325_in = {zll_main_word321_in[31:0], zll_main_word321_in[63:32]};
  assign zll_pure_dispatch110_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word68_in = {zll_pure_dispatch110_in[71:39], zll_pure_dispatch110_in[31:0]};
  assign zll_main_word685_in = {main_word68_in[64:32], main_word68_in[64:32], main_word68_in[31:0]};
  assign zll_main_word683_in = {zll_main_word685_in[97:65], zll_main_word685_in[31:0]};
  assign zll_main_word682_in = {zll_main_word683_in[31:0], zll_main_word683_in[64:32]};
  assign zll_main_word68_in = zll_main_word682_in[64:33];
  assign zll_main_word681_in = {zll_main_word685_in[31:0], zll_main_word685_in[64:32]};
  assign zll_main_word684_in = {zll_main_word681_in[64:33], zll_main_word681_in[31:0]};
  assign zll_main_word686_in = {zll_main_word684_in[31:0], zll_main_word684_in[63:32]};
  assign zll_pure_dispatch93_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word37_in = {zll_pure_dispatch93_in[71:39], zll_pure_dispatch93_in[31:0]};
  assign zll_main_word373_in = {main_word37_in[64:32], main_word37_in[64:32], main_word37_in[31:0]};
  assign zll_main_word377_in = {zll_main_word373_in[97:65], zll_main_word373_in[31:0]};
  assign zll_main_word372_in = {zll_main_word377_in[31:0], zll_main_word377_in[64:32]};
  assign zll_main_word375_in = zll_main_word372_in[64:33];
  assign zll_main_word374_in = {zll_main_word373_in[31:0], zll_main_word373_in[64:32]};
  assign zll_main_word376_in = {zll_main_word374_in[64:33], zll_main_word374_in[31:0]};
  assign zll_main_word371_in = {zll_main_word376_in[31:0], zll_main_word376_in[63:32]};
  assign zll_pure_dispatch58_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word58_in = {zll_pure_dispatch58_in[71:39], zll_pure_dispatch58_in[31:0]};
  assign zll_main_word586_in = {main_word58_in[64:32], main_word58_in[64:32], main_word58_in[31:0]};
  assign zll_main_word583_in = {zll_main_word586_in[97:65], zll_main_word586_in[31:0]};
  assign zll_main_word584_in = {zll_main_word583_in[31:0], zll_main_word583_in[64:32]};
  assign zll_main_word58_in = zll_main_word584_in[64:33];
  assign zll_main_word582_in = {zll_main_word586_in[31:0], zll_main_word586_in[64:32]};
  assign zll_main_word581_in = {zll_main_word582_in[64:33], zll_main_word582_in[31:0]};
  assign zll_main_word585_in = {zll_main_word581_in[31:0], zll_main_word581_in[63:32]};
  assign zll_pure_dispatch92_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word31_in = {zll_pure_dispatch92_in[71:39], zll_pure_dispatch92_in[31:0]};
  assign zll_main_word315_in = {main_word31_in[64:32], main_word31_in[64:32], main_word31_in[31:0]};
  assign zll_main_word311_in = {zll_main_word315_in[97:65], zll_main_word315_in[31:0]};
  assign zll_main_word3110_in = {zll_main_word311_in[31:0], zll_main_word311_in[64:32]};
  assign zll_main_word319_in = zll_main_word3110_in[64:33];
  assign zll_main_word31_in = {zll_main_word315_in[31:0], zll_main_word315_in[64:32]};
  assign zll_main_word312_in = {zll_main_word31_in[64:33], zll_main_word31_in[31:0]};
  assign zll_main_word3111_in = {zll_main_word312_in[31:0], zll_main_word312_in[63:32]};
  assign zll_pure_dispatch15_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word82_in = {zll_pure_dispatch15_in[71:39], zll_pure_dispatch15_in[31:0]};
  assign zll_main_word821_in = {main_word82_in[64:32], main_word82_in[64:32], main_word82_in[31:0]};
  assign zll_main_word823_in = {zll_main_word821_in[97:65], zll_main_word821_in[31:0]};
  assign zll_main_word824_in = {zll_main_word823_in[31:0], zll_main_word823_in[64:32]};
  assign zll_main_word825_in = zll_main_word824_in[64:33];
  assign zll_main_word822_in = {zll_main_word821_in[31:0], zll_main_word821_in[64:32]};
  assign zll_main_word826_in = {zll_main_word822_in[64:33], zll_main_word822_in[31:0]};
  assign zll_main_word827_in = {zll_main_word826_in[31:0], zll_main_word826_in[63:32]};
  assign zll_pure_dispatch86_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word52_in = {zll_pure_dispatch86_in[71:39], zll_pure_dispatch86_in[31:0]};
  assign zll_main_word525_in = {main_word52_in[64:32], main_word52_in[64:32], main_word52_in[31:0]};
  assign zll_main_word524_in = {zll_main_word525_in[97:65], zll_main_word525_in[31:0]};
  assign zll_main_word5210_in = {zll_main_word524_in[31:0], zll_main_word524_in[64:32]};
  assign zll_main_word521_in = zll_main_word5210_in[64:33];
  assign zll_main_word526_in = {zll_main_word525_in[31:0], zll_main_word525_in[64:32]};
  assign zll_main_word522_in = {zll_main_word526_in[64:33], zll_main_word526_in[31:0]};
  assign zll_main_word523_in = {zll_main_word522_in[31:0], zll_main_word522_in[63:32]};
  assign zll_pure_dispatch8_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word101_in = {zll_pure_dispatch8_in[71:39], zll_pure_dispatch8_in[31:0]};
  assign zll_main_word1011_in = {main_word101_in[64:32], main_word101_in[64:32], main_word101_in[31:0]};
  assign zll_main_word1016_in = {zll_main_word1011_in[97:65], zll_main_word1011_in[31:0]};
  assign zll_main_word1019_in = {zll_main_word1016_in[31:0], zll_main_word1016_in[64:32]};
  assign zll_main_word1012_in = zll_main_word1019_in[64:33];
  assign zll_main_word10110_in = {zll_main_word1011_in[31:0], zll_main_word1011_in[64:32]};
  assign zll_main_word1014_in = {zll_main_word10110_in[64:33], zll_main_word10110_in[31:0]};
  assign zll_main_word1013_in = {zll_main_word1014_in[31:0], zll_main_word1014_in[63:32]};
  assign zll_pure_dispatch116_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word80_in = {zll_pure_dispatch116_in[71:39], zll_pure_dispatch116_in[31:0]};
  assign zll_main_word803_in = {main_word80_in[64:32], main_word80_in[64:32], main_word80_in[31:0]};
  assign zll_main_word802_in = {zll_main_word803_in[97:65], zll_main_word803_in[31:0]};
  assign zll_main_word804_in = {zll_main_word802_in[31:0], zll_main_word802_in[64:32]};
  assign zll_main_word801_in = zll_main_word804_in[64:33];
  assign zll_main_word806_in = {zll_main_word803_in[31:0], zll_main_word803_in[64:32]};
  assign zll_main_word80_in = {zll_main_word806_in[64:33], zll_main_word806_in[31:0]};
  assign zll_main_word805_in = {zll_main_word80_in[31:0], zll_main_word80_in[63:32]};
  assign zll_pure_dispatch90_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word39_in = {zll_pure_dispatch90_in[71:39], zll_pure_dispatch90_in[31:0]};
  assign zll_main_word39_in = {main_word39_in[64:32], main_word39_in[64:32], main_word39_in[31:0]};
  assign zll_main_word395_in = {zll_main_word39_in[97:65], zll_main_word39_in[31:0]};
  assign zll_main_word393_in = {zll_main_word395_in[31:0], zll_main_word395_in[64:32]};
  assign zll_main_word391_in = zll_main_word393_in[64:33];
  assign zll_main_word392_in = {zll_main_word39_in[31:0], zll_main_word39_in[64:32]};
  assign zll_main_word394_in = {zll_main_word392_in[64:33], zll_main_word392_in[31:0]};
  assign zll_main_word396_in = {zll_main_word394_in[31:0], zll_main_word394_in[63:32]};
  assign zll_pure_dispatch7_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word21_in = {zll_pure_dispatch7_in[71:39], zll_pure_dispatch7_in[31:0]};
  assign zll_main_word216_in = {main_word21_in[64:32], main_word21_in[64:32], main_word21_in[31:0]};
  assign zll_main_word2110_in = {zll_main_word216_in[97:65], zll_main_word216_in[31:0]};
  assign zll_main_word2112_in = {zll_main_word2110_in[31:0], zll_main_word2110_in[64:32]};
  assign zll_main_word218_in = zll_main_word2112_in[64:33];
  assign zll_main_word2111_in = {zll_main_word216_in[31:0], zll_main_word216_in[64:32]};
  assign zll_main_word217_in = {zll_main_word2111_in[64:33], zll_main_word2111_in[31:0]};
  assign zll_main_word2113_in = {zll_main_word217_in[31:0], zll_main_word217_in[63:32]};
  assign zll_pure_dispatch88_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word16_in = {zll_pure_dispatch88_in[71:39], zll_pure_dispatch88_in[31:0]};
  assign zll_main_word164_in = {main_word16_in[64:32], main_word16_in[64:32], main_word16_in[31:0]};
  assign zll_main_word163_in = {zll_main_word164_in[97:65], zll_main_word164_in[31:0]};
  assign zll_main_word162_in = {zll_main_word163_in[31:0], zll_main_word163_in[64:32]};
  assign zll_main_word165_in = zll_main_word162_in[64:33];
  assign zll_main_word161_in = {zll_main_word164_in[31:0], zll_main_word164_in[64:32]};
  assign zll_main_word166_in = {zll_main_word161_in[64:33], zll_main_word161_in[31:0]};
  assign zll_main_word16_in = {zll_main_word166_in[31:0], zll_main_word166_in[63:32]};
  assign zll_pure_dispatch97_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word112_in = {zll_pure_dispatch97_in[71:39], zll_pure_dispatch97_in[31:0]};
  assign zll_main_word112_in = {main_word112_in[64:32], main_word112_in[64:32], main_word112_in[31:0]};
  assign zll_main_word1121_in = {zll_main_word112_in[97:65], zll_main_word112_in[31:0]};
  assign zll_main_word1123_in = {zll_main_word1121_in[31:0], zll_main_word1121_in[64:32]};
  assign zll_main_word1126_in = zll_main_word1123_in[64:33];
  assign zll_main_word1122_in = {zll_main_word112_in[31:0], zll_main_word112_in[64:32]};
  assign zll_main_word1124_in = {zll_main_word1122_in[64:33], zll_main_word1122_in[31:0]};
  assign zll_main_word1125_in = {zll_main_word1124_in[31:0], zll_main_word1124_in[63:32]};
  assign zll_pure_dispatch80_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word12_in = {zll_pure_dispatch80_in[71:39], zll_pure_dispatch80_in[31:0]};
  assign zll_main_word124_in = {main_word12_in[64:32], main_word12_in[64:32], main_word12_in[31:0]};
  assign zll_main_word1215_in = {zll_main_word124_in[97:65], zll_main_word124_in[31:0]};
  assign zll_main_word1219_in = {zll_main_word1215_in[31:0], zll_main_word1215_in[64:32]};
  assign zll_main_word1210_in = zll_main_word1219_in[64:33];
  assign zll_main_word127_in = {zll_main_word124_in[31:0], zll_main_word124_in[64:32]};
  assign zll_main_word1211_in = {zll_main_word127_in[64:33], zll_main_word127_in[31:0]};
  assign zll_main_word1213_in = {zll_main_word1211_in[31:0], zll_main_word1211_in[63:32]};
  assign zll_pure_dispatch87_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word42_in = {zll_pure_dispatch87_in[71:39], zll_pure_dispatch87_in[31:0]};
  assign zll_main_word429_in = {main_word42_in[64:32], main_word42_in[64:32], main_word42_in[31:0]};
  assign zll_main_word421_in = {zll_main_word429_in[97:65], zll_main_word429_in[31:0]};
  assign zll_main_word4210_in = {zll_main_word421_in[31:0], zll_main_word421_in[64:32]};
  assign zll_main_word4212_in = zll_main_word4210_in[64:33];
  assign zll_main_word42_in = {zll_main_word429_in[31:0], zll_main_word429_in[64:32]};
  assign zll_main_word4211_in = {zll_main_word42_in[64:33], zll_main_word42_in[31:0]};
  assign zll_main_word424_in = {zll_main_word4211_in[31:0], zll_main_word4211_in[63:32]};
  assign zll_pure_dispatch57_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word1_in = {zll_pure_dispatch57_in[71:39], zll_pure_dispatch57_in[31:0]};
  assign zll_main_word121_in = {main_word1_in[64:32], main_word1_in[64:32], main_word1_in[31:0]};
  assign zll_main_word147_in = {zll_main_word121_in[97:65], zll_main_word121_in[31:0]};
  assign zll_main_word09_in = {zll_main_word147_in[31:0], zll_main_word147_in[64:32]};
  ZLL_Main_word09  instR2 (zll_main_word09_in[64:33], zll_main_word09_out);
  assign zll_main_word130_in = {zll_main_word121_in[31:0], zll_main_word121_in[64:32]};
  assign zll_main_word138_in = {zll_main_word130_in[64:33], zll_main_word130_in[31:0]};
  assign zll_main_word133_in = {zll_main_word138_in[31:0], zll_main_word138_in[63:32]};
  assign zll_main_word430_inR1 = {zll_main_word133_in[31:0], zll_main_word133_in[31:0]};
  ZLL_Main_word430  instR3 (zll_main_word430_inR1[63:0], zll_main_word430_outR1);
  assign zll_main_word12_in = {zll_main_word133_in[63:32], zll_main_word430_outR1};
  assign zll_main_word140_in = {zll_main_word12_in[97:66], zll_main_word12_in[65:0]};
  assign zll_main_word128_in = {zll_main_word140_in[97:66], zll_main_word140_in[63:32], zll_main_word140_in[31:0]};
  assign test1_in = {zll_main_word128_in[95:64], zll_main_word128_in[63:32]};
  test1  instR4 (test1_in[63:32], test1_in[31:0], extresR1[0]);
  assign zll_pure_dispatch111_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word41_in = {zll_pure_dispatch111_in[71:39], zll_pure_dispatch111_in[31:0]};
  assign zll_main_word413_in = {main_word41_in[64:32], main_word41_in[64:32], main_word41_in[31:0]};
  assign zll_main_word411_in = {zll_main_word413_in[97:65], zll_main_word413_in[31:0]};
  assign zll_main_word415_in = {zll_main_word411_in[31:0], zll_main_word411_in[64:32]};
  assign zll_main_word416_in = zll_main_word415_in[64:33];
  assign zll_main_word414_in = {zll_main_word413_in[31:0], zll_main_word413_in[64:32]};
  assign zll_main_word4110_in = {zll_main_word414_in[64:33], zll_main_word414_in[31:0]};
  assign zll_main_word412_in = {zll_main_word4110_in[31:0], zll_main_word4110_in[63:32]};
  assign zll_pure_dispatch32_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word96_in = {zll_pure_dispatch32_in[71:39], zll_pure_dispatch32_in[31:0]};
  assign zll_main_word966_in = {main_word96_in[64:32], main_word96_in[64:32], main_word96_in[31:0]};
  assign zll_main_word961_in = {zll_main_word966_in[97:65], zll_main_word966_in[31:0]};
  assign zll_main_word964_in = {zll_main_word961_in[31:0], zll_main_word961_in[64:32]};
  assign zll_main_word963_in = zll_main_word964_in[64:33];
  assign zll_main_word965_in = {zll_main_word966_in[31:0], zll_main_word966_in[64:32]};
  assign zll_main_word96_in = {zll_main_word965_in[64:33], zll_main_word965_in[31:0]};
  assign zll_main_word962_in = {zll_main_word96_in[31:0], zll_main_word96_in[63:32]};
  assign zll_pure_dispatch79_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word53_in = {zll_pure_dispatch79_in[71:39], zll_pure_dispatch79_in[31:0]};
  assign zll_main_word535_in = {main_word53_in[64:32], main_word53_in[64:32], main_word53_in[31:0]};
  assign zll_main_word53_in = {zll_main_word535_in[97:65], zll_main_word535_in[31:0]};
  assign zll_main_word532_in = {zll_main_word53_in[31:0], zll_main_word53_in[64:32]};
  assign zll_main_word533_in = zll_main_word532_in[64:33];
  assign zll_main_word531_in = {zll_main_word535_in[31:0], zll_main_word535_in[64:32]};
  assign zll_main_word536_in = {zll_main_word531_in[64:33], zll_main_word531_in[31:0]};
  assign zll_main_word534_in = {zll_main_word536_in[31:0], zll_main_word536_in[63:32]};
  assign zll_pure_dispatch44_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word89_in = {zll_pure_dispatch44_in[71:39], zll_pure_dispatch44_in[31:0]};
  assign zll_main_word894_in = {main_word89_in[64:32], main_word89_in[64:32], main_word89_in[31:0]};
  assign zll_main_word896_in = {zll_main_word894_in[97:65], zll_main_word894_in[31:0]};
  assign zll_main_word892_in = {zll_main_word896_in[31:0], zll_main_word896_in[64:32]};
  assign zll_main_word895_in = zll_main_word892_in[64:33];
  assign zll_main_word891_in = {zll_main_word894_in[31:0], zll_main_word894_in[64:32]};
  assign zll_main_word89_in = {zll_main_word891_in[64:33], zll_main_word891_in[31:0]};
  assign zll_main_word893_in = {zll_main_word89_in[31:0], zll_main_word89_in[63:32]};
  assign zll_pure_dispatch82_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word35_in = {zll_pure_dispatch82_in[71:39], zll_pure_dispatch82_in[31:0]};
  assign zll_main_word353_in = {main_word35_in[64:32], main_word35_in[64:32], main_word35_in[31:0]};
  assign zll_main_word35_in = {zll_main_word353_in[97:65], zll_main_word353_in[31:0]};
  assign zll_main_word351_in = {zll_main_word35_in[31:0], zll_main_word35_in[64:32]};
  assign zll_main_word354_in = zll_main_word351_in[64:33];
  assign zll_main_word352_in = {zll_main_word353_in[31:0], zll_main_word353_in[64:32]};
  assign zll_main_word355_in = {zll_main_word352_in[64:33], zll_main_word352_in[31:0]};
  assign zll_main_word356_in = {zll_main_word355_in[31:0], zll_main_word355_in[63:32]};
  assign zll_pure_dispatch19_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word94_in = {zll_pure_dispatch19_in[71:39], zll_pure_dispatch19_in[31:0]};
  assign zll_main_word94_in = {main_word94_in[64:32], main_word94_in[64:32], main_word94_in[31:0]};
  assign zll_main_word945_in = {zll_main_word94_in[97:65], zll_main_word94_in[31:0]};
  assign zll_main_word944_in = {zll_main_word945_in[31:0], zll_main_word945_in[64:32]};
  assign zll_main_word946_in = zll_main_word944_in[64:33];
  assign zll_main_word943_in = {zll_main_word94_in[31:0], zll_main_word94_in[64:32]};
  assign zll_main_word942_in = {zll_main_word943_in[64:33], zll_main_word943_in[31:0]};
  assign zll_main_word941_in = {zll_main_word942_in[31:0], zll_main_word942_in[63:32]};
  assign zll_pure_dispatch71_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word55_in = {zll_pure_dispatch71_in[71:39], zll_pure_dispatch71_in[31:0]};
  assign zll_main_word55_in = {main_word55_in[64:32], main_word55_in[64:32], main_word55_in[31:0]};
  assign zll_main_word552_in = {zll_main_word55_in[97:65], zll_main_word55_in[31:0]};
  assign zll_main_word551_in = {zll_main_word552_in[31:0], zll_main_word552_in[64:32]};
  assign zll_main_word556_in = zll_main_word551_in[64:33];
  assign zll_main_word553_in = {zll_main_word55_in[31:0], zll_main_word55_in[64:32]};
  assign zll_main_word555_in = {zll_main_word553_in[64:33], zll_main_word553_in[31:0]};
  assign zll_main_word554_in = {zll_main_word555_in[31:0], zll_main_word555_in[63:32]};
  assign zll_pure_dispatch48_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word26_in = {zll_pure_dispatch48_in[71:39], zll_pure_dispatch48_in[31:0]};
  assign zll_main_word266_in = {main_word26_in[64:32], main_word26_in[64:32], main_word26_in[31:0]};
  assign zll_main_word264_in = {zll_main_word266_in[97:65], zll_main_word266_in[31:0]};
  assign zll_main_word263_in = {zll_main_word264_in[31:0], zll_main_word264_in[64:32]};
  assign zll_main_word261_in = zll_main_word263_in[64:33];
  assign zll_main_word26_in = {zll_main_word266_in[31:0], zll_main_word266_in[64:32]};
  assign zll_main_word265_in = {zll_main_word26_in[64:33], zll_main_word26_in[31:0]};
  assign zll_main_word262_in = {zll_main_word265_in[31:0], zll_main_word265_in[63:32]};
  assign zll_pure_dispatch77_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word123_in = {zll_pure_dispatch77_in[71:39], zll_pure_dispatch77_in[31:0]};
  assign zll_main_word1236_in = {main_word123_in[64:32], main_word123_in[64:32], main_word123_in[31:0]};
  assign zll_main_word1231_in = {zll_main_word1236_in[97:65], zll_main_word1236_in[31:0]};
  assign zll_main_word1233_in = {zll_main_word1231_in[31:0], zll_main_word1231_in[64:32]};
  assign zll_main_word1235_in = zll_main_word1233_in[64:33];
  assign zll_main_word1232_in = {zll_main_word1236_in[31:0], zll_main_word1236_in[64:32]};
  assign zll_main_word123_in = {zll_main_word1232_in[64:33], zll_main_word1232_in[31:0]};
  assign zll_main_word1234_in = {zll_main_word123_in[31:0], zll_main_word123_in[63:32]};
  assign zll_pure_dispatch27_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word27_in = {zll_pure_dispatch27_in[71:39], zll_pure_dispatch27_in[31:0]};
  assign zll_main_word271_in = {main_word27_in[64:32], main_word27_in[64:32], main_word27_in[31:0]};
  assign zll_main_word272_in = {zll_main_word271_in[97:65], zll_main_word271_in[31:0]};
  assign zll_main_word27_in = {zll_main_word272_in[31:0], zll_main_word272_in[64:32]};
  assign zll_main_word273_in = zll_main_word27_in[64:33];
  assign zll_main_word275_in = {zll_main_word271_in[31:0], zll_main_word271_in[64:32]};
  assign zll_main_word274_in = {zll_main_word275_in[64:33], zll_main_word275_in[31:0]};
  assign zll_main_word276_in = {zll_main_word274_in[31:0], zll_main_word274_in[63:32]};
  assign zll_pure_dispatch41_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word83_in = {zll_pure_dispatch41_in[71:39], zll_pure_dispatch41_in[31:0]};
  assign zll_main_word831_in = {main_word83_in[64:32], main_word83_in[64:32], main_word83_in[31:0]};
  assign zll_main_word835_in = {zll_main_word831_in[97:65], zll_main_word831_in[31:0]};
  assign zll_main_word83_in = {zll_main_word835_in[31:0], zll_main_word835_in[64:32]};
  assign zll_main_word833_in = zll_main_word83_in[64:33];
  assign zll_main_word836_in = {zll_main_word831_in[31:0], zll_main_word831_in[64:32]};
  assign zll_main_word832_in = {zll_main_word836_in[64:33], zll_main_word836_in[31:0]};
  assign zll_main_word834_in = {zll_main_word832_in[31:0], zll_main_word832_in[63:32]};
  assign zll_pure_dispatch117_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word13_in = {zll_pure_dispatch117_in[71:39], zll_pure_dispatch117_in[31:0]};
  assign zll_main_word137_in = {main_word13_in[64:32], main_word13_in[64:32], main_word13_in[31:0]};
  assign zll_main_word132_in = {zll_main_word137_in[97:65], zll_main_word137_in[31:0]};
  assign zll_main_word131_in = {zll_main_word132_in[31:0], zll_main_word132_in[64:32]};
  assign zll_main_word134_in = zll_main_word131_in[64:33];
  assign zll_main_word13_in = {zll_main_word137_in[31:0], zll_main_word137_in[64:32]};
  assign zll_main_word1311_in = {zll_main_word13_in[64:33], zll_main_word13_in[31:0]};
  assign zll_main_word1310_in = {zll_main_word1311_in[31:0], zll_main_word1311_in[63:32]};
  assign zll_pure_dispatch64_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word69_in = {zll_pure_dispatch64_in[71:39], zll_pure_dispatch64_in[31:0]};
  assign zll_main_word695_in = {main_word69_in[64:32], main_word69_in[64:32], main_word69_in[31:0]};
  assign zll_main_word69_in = {zll_main_word695_in[97:65], zll_main_word695_in[31:0]};
  assign zll_main_word691_in = {zll_main_word69_in[31:0], zll_main_word69_in[64:32]};
  assign zll_main_word693_in = zll_main_word691_in[64:33];
  assign zll_main_word692_in = {zll_main_word695_in[31:0], zll_main_word695_in[64:32]};
  assign zll_main_word696_in = {zll_main_word692_in[64:33], zll_main_word692_in[31:0]};
  assign zll_main_word694_in = {zll_main_word696_in[31:0], zll_main_word696_in[63:32]};
  assign zll_pure_dispatch69_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word115_in = {zll_pure_dispatch69_in[71:39], zll_pure_dispatch69_in[31:0]};
  assign zll_main_word1155_in = {main_word115_in[64:32], main_word115_in[64:32], main_word115_in[31:0]};
  assign zll_main_word1152_in = {zll_main_word1155_in[97:65], zll_main_word1155_in[31:0]};
  assign zll_main_word1153_in = {zll_main_word1152_in[31:0], zll_main_word1152_in[64:32]};
  assign zll_main_word1154_in = zll_main_word1153_in[64:33];
  assign zll_main_word1151_in = {zll_main_word1155_in[31:0], zll_main_word1155_in[64:32]};
  assign zll_main_word115_in = {zll_main_word1151_in[64:33], zll_main_word1151_in[31:0]};
  assign zll_main_word1156_in = {zll_main_word115_in[31:0], zll_main_word115_in[63:32]};
  assign zll_pure_dispatch21_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word87_in = {zll_pure_dispatch21_in[71:39], zll_pure_dispatch21_in[31:0]};
  assign zll_main_word875_in = {main_word87_in[64:32], main_word87_in[64:32], main_word87_in[31:0]};
  assign zll_main_word873_in = {zll_main_word875_in[97:65], zll_main_word875_in[31:0]};
  assign zll_main_word87_in = {zll_main_word873_in[31:0], zll_main_word873_in[64:32]};
  assign zll_main_word874_in = zll_main_word87_in[64:33];
  assign zll_main_word872_in = {zll_main_word875_in[31:0], zll_main_word875_in[64:32]};
  assign zll_main_word871_in = {zll_main_word872_in[64:33], zll_main_word872_in[31:0]};
  assign zll_main_word876_in = {zll_main_word871_in[31:0], zll_main_word871_in[63:32]};
  assign zll_pure_dispatch72_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word25_in = {zll_pure_dispatch72_in[71:39], zll_pure_dispatch72_in[31:0]};
  assign zll_main_word254_in = {main_word25_in[64:32], main_word25_in[64:32], main_word25_in[31:0]};
  assign zll_main_word256_in = {zll_main_word254_in[97:65], zll_main_word254_in[31:0]};
  assign zll_main_word251_in = {zll_main_word256_in[31:0], zll_main_word256_in[64:32]};
  assign zll_main_word252_in = zll_main_word251_in[64:33];
  assign zll_main_word25_in = {zll_main_word254_in[31:0], zll_main_word254_in[64:32]};
  assign zll_main_word253_in = {zll_main_word25_in[64:33], zll_main_word25_in[31:0]};
  assign zll_main_word255_in = {zll_main_word253_in[31:0], zll_main_word253_in[63:32]};
  assign zll_pure_dispatch103_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word19_in = {zll_pure_dispatch103_in[71:39], zll_pure_dispatch103_in[31:0]};
  assign zll_main_word196_in = {main_word19_in[64:32], main_word19_in[64:32], main_word19_in[31:0]};
  assign zll_main_word194_in = {zll_main_word196_in[97:65], zll_main_word196_in[31:0]};
  assign zll_main_word193_in = {zll_main_word194_in[31:0], zll_main_word194_in[64:32]};
  assign zll_main_word19_in = zll_main_word193_in[64:33];
  assign zll_main_word195_in = {zll_main_word196_in[31:0], zll_main_word196_in[64:32]};
  assign zll_main_word191_in = {zll_main_word195_in[64:33], zll_main_word195_in[31:0]};
  assign zll_main_word192_in = {zll_main_word191_in[31:0], zll_main_word191_in[63:32]};
  assign zll_pure_dispatch62_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word76_in = {zll_pure_dispatch62_in[71:39], zll_pure_dispatch62_in[31:0]};
  assign zll_main_word762_in = {main_word76_in[64:32], main_word76_in[64:32], main_word76_in[31:0]};
  assign zll_main_word765_in = {zll_main_word762_in[97:65], zll_main_word762_in[31:0]};
  assign zll_main_word761_in = {zll_main_word765_in[31:0], zll_main_word765_in[64:32]};
  assign zll_main_word763_in = zll_main_word761_in[64:33];
  assign zll_main_word764_in = {zll_main_word762_in[31:0], zll_main_word762_in[64:32]};
  assign zll_main_word767_in = {zll_main_word764_in[64:33], zll_main_word764_in[31:0]};
  assign zll_main_word766_in = {zll_main_word767_in[31:0], zll_main_word767_in[63:32]};
  assign zll_pure_dispatch91_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word85_in = {zll_pure_dispatch91_in[71:39], zll_pure_dispatch91_in[31:0]};
  assign zll_main_word854_in = {main_word85_in[64:32], main_word85_in[64:32], main_word85_in[31:0]};
  assign zll_main_word852_in = {zll_main_word854_in[97:65], zll_main_word854_in[31:0]};
  assign zll_main_word85_in = {zll_main_word852_in[31:0], zll_main_word852_in[64:32]};
  assign zll_main_word856_in = zll_main_word85_in[64:33];
  assign zll_main_word855_in = {zll_main_word854_in[31:0], zll_main_word854_in[64:32]};
  assign zll_main_word853_in = {zll_main_word855_in[64:33], zll_main_word855_in[31:0]};
  assign zll_main_word851_in = {zll_main_word853_in[31:0], zll_main_word853_in[63:32]};
  assign zll_pure_dispatch122_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word91_in = {zll_pure_dispatch122_in[71:39], zll_pure_dispatch122_in[31:0]};
  assign zll_main_word91_in = {main_word91_in[64:32], main_word91_in[64:32], main_word91_in[31:0]};
  assign zll_main_word913_in = {zll_main_word91_in[97:65], zll_main_word91_in[31:0]};
  assign zll_main_word912_in = {zll_main_word913_in[31:0], zll_main_word913_in[64:32]};
  assign zll_main_word915_in = zll_main_word912_in[64:33];
  assign zll_main_word911_in = {zll_main_word91_in[31:0], zll_main_word91_in[64:32]};
  assign zll_main_word914_in = {zll_main_word911_in[64:33], zll_main_word911_in[31:0]};
  assign zll_main_word916_in = {zll_main_word914_in[31:0], zll_main_word914_in[63:32]};
  assign zll_pure_dispatch13_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word5_in = {zll_pure_dispatch13_in[71:39], zll_pure_dispatch13_in[31:0]};
  assign zll_main_word515_in = {main_word5_in[64:32], main_word5_in[64:32], main_word5_in[31:0]};
  assign zll_main_word527_in = {zll_main_word515_in[97:65], zll_main_word515_in[31:0]};
  assign zll_main_word519_in = {zll_main_word527_in[31:0], zll_main_word527_in[64:32]};
  assign zll_main_word517_in = zll_main_word519_in[64:33];
  assign zll_main_word528_in = {zll_main_word515_in[31:0], zll_main_word515_in[64:32]};
  assign zll_main_word54_in = {zll_main_word528_in[64:33], zll_main_word528_in[31:0]};
  assign zll_main_word513_in = {zll_main_word54_in[31:0], zll_main_word54_in[63:32]};
  assign zll_main_word430_inR2 = {zll_main_word513_in[31:0], zll_main_word513_in[31:0]};
  ZLL_Main_word430  instR5 (zll_main_word430_inR2[63:0], zll_main_word430_outR2);
  assign zll_main_word5_in = {zll_main_word513_in[63:32], zll_main_word430_outR2};
  assign zll_main_word530_in = {zll_main_word5_in[97:66], zll_main_word5_in[65:0]};
  assign zll_main_word514_in = {zll_main_word530_in[97:66], zll_main_word530_in[63:32], zll_main_word530_in[31:0]};
  assign test3_in = {zll_main_word514_in[95:64], zll_main_word514_in[63:32]};
  test3  instR6 (test3_in[63:32], test3_in[31:0], extresR2[0]);
  assign zll_pure_dispatch6_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word75_in = {zll_pure_dispatch6_in[71:39], zll_pure_dispatch6_in[31:0]};
  assign zll_main_word755_in = {main_word75_in[64:32], main_word75_in[64:32], main_word75_in[31:0]};
  assign zll_main_word756_in = {zll_main_word755_in[97:65], zll_main_word755_in[31:0]};
  assign zll_main_word754_in = {zll_main_word756_in[31:0], zll_main_word756_in[64:32]};
  assign zll_main_word75_in = zll_main_word754_in[64:33];
  assign zll_main_word753_in = {zll_main_word755_in[31:0], zll_main_word755_in[64:32]};
  assign zll_main_word752_in = {zll_main_word753_in[64:33], zll_main_word753_in[31:0]};
  assign zll_main_word751_in = {zll_main_word752_in[31:0], zll_main_word752_in[63:32]};
  assign zll_pure_dispatch66_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word86_in = {zll_pure_dispatch66_in[71:39], zll_pure_dispatch66_in[31:0]};
  assign zll_main_word862_in = {main_word86_in[64:32], main_word86_in[64:32], main_word86_in[31:0]};
  assign zll_main_word861_in = {zll_main_word862_in[97:65], zll_main_word862_in[31:0]};
  assign zll_main_word865_in = {zll_main_word861_in[31:0], zll_main_word861_in[64:32]};
  assign zll_main_word864_in = zll_main_word865_in[64:33];
  assign zll_main_word86_in = {zll_main_word862_in[31:0], zll_main_word862_in[64:32]};
  assign zll_main_word866_in = {zll_main_word86_in[64:33], zll_main_word86_in[31:0]};
  assign zll_main_word863_in = {zll_main_word866_in[31:0], zll_main_word866_in[63:32]};
  assign zll_pure_dispatch17_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word7_in = {zll_pure_dispatch17_in[71:39], zll_pure_dispatch17_in[31:0]};
  assign zll_main_word7_in = {main_word7_in[64:32], main_word7_in[64:32], main_word7_in[31:0]};
  assign zll_main_word717_in = {zll_main_word7_in[97:65], zll_main_word7_in[31:0]};
  assign zll_main_word720_in = {zll_main_word717_in[31:0], zll_main_word717_in[64:32]};
  assign zll_main_word715_in = zll_main_word720_in[64:33];
  assign zll_main_word710_in = {zll_main_word7_in[31:0], zll_main_word7_in[64:32]};
  assign zll_main_word76_in = {zll_main_word710_in[64:33], zll_main_word710_in[31:0]};
  assign zll_main_word714_in = {zll_main_word76_in[31:0], zll_main_word76_in[63:32]};
  assign zll_pure_dispatch63_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word3_in = {zll_pure_dispatch63_in[71:39], zll_pure_dispatch63_in[31:0]};
  assign zll_main_word337_in = {main_word3_in[64:32], main_word3_in[64:32], main_word3_in[31:0]};
  assign zll_main_word310_in = {zll_main_word337_in[97:65], zll_main_word337_in[31:0]};
  assign zll_main_word314_in = {zll_main_word310_in[31:0], zll_main_word310_in[64:32]};
  ZLL_Main_word314  instR7 (zll_main_word314_in[64:33], zll_main_word314_out);
  assign zll_main_word37_in = {zll_main_word337_in[31:0], zll_main_word337_in[64:32]};
  assign zll_main_word313_in = {zll_main_word37_in[64:33], zll_main_word37_in[31:0]};
  assign zll_main_word317_in = {zll_main_word313_in[31:0], zll_main_word313_in[63:32]};
  assign zll_main_word430_inR3 = {zll_main_word317_in[31:0], zll_main_word317_in[31:0]};
  ZLL_Main_word430  instR8 (zll_main_word430_inR3[63:0], zll_main_word430_outR3);
  assign zll_main_word33_in = {zll_main_word317_in[63:32], zll_main_word430_outR3};
  assign zll_main_word329_in = {zll_main_word33_in[97:66], zll_main_word33_in[65:0]};
  assign zll_main_word3_in = {zll_main_word329_in[97:66], zll_main_word329_in[63:32], zll_main_word329_in[31:0]};
  assign test1_inR1 = {zll_main_word3_in[95:64], zll_main_word3_in[63:32]};
  test1  instR9 (test1_inR1[63:32], test1_inR1[31:0], extresR3[0]);
  assign zll_pure_dispatch112_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word45_in = {zll_pure_dispatch112_in[71:39], zll_pure_dispatch112_in[31:0]};
  assign zll_main_word456_in = {main_word45_in[64:32], main_word45_in[64:32], main_word45_in[31:0]};
  assign zll_main_word45_in = {zll_main_word456_in[97:65], zll_main_word456_in[31:0]};
  assign zll_main_word455_in = {zll_main_word45_in[31:0], zll_main_word45_in[64:32]};
  assign zll_main_word453_in = zll_main_word455_in[64:33];
  assign zll_main_word451_in = {zll_main_word456_in[31:0], zll_main_word456_in[64:32]};
  assign zll_main_word452_in = {zll_main_word451_in[64:33], zll_main_word451_in[31:0]};
  assign zll_main_word454_in = {zll_main_word452_in[31:0], zll_main_word452_in[63:32]};
  assign zll_pure_dispatch26_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word43_in = {zll_pure_dispatch26_in[71:39], zll_pure_dispatch26_in[31:0]};
  assign zll_main_word433_in = {main_word43_in[64:32], main_word43_in[64:32], main_word43_in[31:0]};
  assign zll_main_word435_in = {zll_main_word433_in[97:65], zll_main_word433_in[31:0]};
  assign zll_main_word437_in = {zll_main_word435_in[31:0], zll_main_word435_in[64:32]};
  assign zll_main_word432_in = zll_main_word437_in[64:33];
  assign zll_main_word431_in = {zll_main_word433_in[31:0], zll_main_word433_in[64:32]};
  assign zll_main_word434_in = {zll_main_word431_in[64:33], zll_main_word431_in[31:0]};
  assign zll_main_word436_in = {zll_main_word434_in[31:0], zll_main_word434_in[63:32]};
  assign zll_pure_dispatch_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word116_in = {zll_pure_dispatch_in[71:39], zll_pure_dispatch_in[31:0]};
  assign zll_main_word1166_in = {main_word116_in[64:32], main_word116_in[64:32], main_word116_in[31:0]};
  assign zll_main_word1167_in = {zll_main_word1166_in[97:65], zll_main_word1166_in[31:0]};
  assign zll_main_word1165_in = {zll_main_word1167_in[31:0], zll_main_word1167_in[64:32]};
  assign zll_main_word1162_in = zll_main_word1165_in[64:33];
  assign zll_main_word1161_in = {zll_main_word1166_in[31:0], zll_main_word1166_in[64:32]};
  assign zll_main_word1164_in = {zll_main_word1161_in[64:33], zll_main_word1161_in[31:0]};
  assign zll_main_word1163_in = {zll_main_word1164_in[31:0], zll_main_word1164_in[63:32]};
  assign zll_pure_dispatch118_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word54_in = {zll_pure_dispatch118_in[71:39], zll_pure_dispatch118_in[31:0]};
  assign zll_main_word541_in = {main_word54_in[64:32], main_word54_in[64:32], main_word54_in[31:0]};
  assign zll_main_word547_in = {zll_main_word541_in[97:65], zll_main_word541_in[31:0]};
  assign zll_main_word543_in = {zll_main_word547_in[31:0], zll_main_word547_in[64:32]};
  assign zll_main_word542_in = zll_main_word543_in[64:33];
  assign zll_main_word545_in = {zll_main_word541_in[31:0], zll_main_word541_in[64:32]};
  assign zll_main_word546_in = {zll_main_word545_in[64:33], zll_main_word545_in[31:0]};
  assign zll_main_word544_in = {zll_main_word546_in[31:0], zll_main_word546_in[63:32]};
  assign zll_pure_dispatch126_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word113_in = {zll_pure_dispatch126_in[71:39], zll_pure_dispatch126_in[31:0]};
  assign zll_main_word1135_in = {main_word113_in[64:32], main_word113_in[64:32], main_word113_in[31:0]};
  assign zll_main_word1134_in = {zll_main_word1135_in[97:65], zll_main_word1135_in[31:0]};
  assign zll_main_word1136_in = {zll_main_word1134_in[31:0], zll_main_word1134_in[64:32]};
  assign zll_main_word1132_in = zll_main_word1136_in[64:33];
  assign zll_main_word1131_in = {zll_main_word1135_in[31:0], zll_main_word1135_in[64:32]};
  assign zll_main_word1133_in = {zll_main_word1131_in[64:33], zll_main_word1131_in[31:0]};
  assign zll_main_word113_in = {zll_main_word1133_in[31:0], zll_main_word1133_in[63:32]};
  assign zll_pure_dispatch83_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word47_in = {zll_pure_dispatch83_in[71:39], zll_pure_dispatch83_in[31:0]};
  assign zll_main_word474_in = {main_word47_in[64:32], main_word47_in[64:32], main_word47_in[31:0]};
  assign zll_main_word471_in = {zll_main_word474_in[97:65], zll_main_word474_in[31:0]};
  assign zll_main_word473_in = {zll_main_word471_in[31:0], zll_main_word471_in[64:32]};
  assign zll_main_word47_in = zll_main_word473_in[64:33];
  assign zll_main_word476_in = {zll_main_word474_in[31:0], zll_main_word474_in[64:32]};
  assign zll_main_word472_in = {zll_main_word476_in[64:33], zll_main_word476_in[31:0]};
  assign zll_main_word475_in = {zll_main_word472_in[31:0], zll_main_word472_in[63:32]};
  assign zll_pure_dispatch102_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word60_in = {zll_pure_dispatch102_in[71:39], zll_pure_dispatch102_in[31:0]};
  assign zll_main_word606_in = {main_word60_in[64:32], main_word60_in[64:32], main_word60_in[31:0]};
  assign zll_main_word60_in = {zll_main_word606_in[97:65], zll_main_word606_in[31:0]};
  assign zll_main_word603_in = {zll_main_word60_in[31:0], zll_main_word60_in[64:32]};
  assign zll_main_word604_in = zll_main_word603_in[64:33];
  assign zll_main_word605_in = {zll_main_word606_in[31:0], zll_main_word606_in[64:32]};
  assign zll_main_word602_in = {zll_main_word605_in[64:33], zll_main_word605_in[31:0]};
  assign zll_main_word601_in = {zll_main_word602_in[31:0], zll_main_word602_in[63:32]};
  assign zll_pure_dispatch33_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word72_in = {zll_pure_dispatch33_in[71:39], zll_pure_dispatch33_in[31:0]};
  assign zll_main_word725_in = {main_word72_in[64:32], main_word72_in[64:32], main_word72_in[31:0]};
  assign zll_main_word72_in = {zll_main_word725_in[97:65], zll_main_word725_in[31:0]};
  assign zll_main_word721_in = {zll_main_word72_in[31:0], zll_main_word72_in[64:32]};
  assign zll_main_word723_in = zll_main_word721_in[64:33];
  assign zll_main_word722_in = {zll_main_word725_in[31:0], zll_main_word725_in[64:32]};
  assign zll_main_word726_in = {zll_main_word722_in[64:33], zll_main_word722_in[31:0]};
  assign zll_main_word724_in = {zll_main_word726_in[31:0], zll_main_word726_in[63:32]};
  assign zll_pure_dispatch50_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word79_in = {zll_pure_dispatch50_in[71:39], zll_pure_dispatch50_in[31:0]};
  assign zll_main_word791_in = {main_word79_in[64:32], main_word79_in[64:32], main_word79_in[31:0]};
  assign zll_main_word796_in = {zll_main_word791_in[97:65], zll_main_word791_in[31:0]};
  assign zll_main_word79_in = {zll_main_word796_in[31:0], zll_main_word796_in[64:32]};
  assign zll_main_word795_in = zll_main_word79_in[64:33];
  assign zll_main_word794_in = {zll_main_word791_in[31:0], zll_main_word791_in[64:32]};
  assign zll_main_word793_in = {zll_main_word794_in[64:33], zll_main_word794_in[31:0]};
  assign zll_main_word792_in = {zll_main_word793_in[31:0], zll_main_word793_in[63:32]};
  assign zll_pure_dispatch56_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word6_in = {zll_pure_dispatch56_in[71:39], zll_pure_dispatch56_in[31:0]};
  assign zll_main_word65_in = {main_word6_in[64:32], main_word6_in[64:32], main_word6_in[31:0]};
  assign zll_main_word629_in = {zll_main_word65_in[97:65], zll_main_word65_in[31:0]};
  assign zll_main_word610_in = {zll_main_word629_in[31:0], zll_main_word629_in[64:32]};
  assign zll_main_word611_in = zll_main_word610_in[64:33];
  assign zll_main_word617_in = {zll_main_word65_in[31:0], zll_main_word65_in[64:32]};
  assign zll_main_word619_in = {zll_main_word617_in[64:33], zll_main_word617_in[31:0]};
  assign zll_main_word6_in = {zll_main_word619_in[31:0], zll_main_word619_in[63:32]};
  assign zll_main_word430_inR4 = {zll_main_word6_in[31:0], zll_main_word6_in[31:0]};
  ZLL_Main_word430  instR10 (zll_main_word430_inR4[63:0], zll_main_word430_outR4);
  assign zll_main_word626_in = {zll_main_word6_in[63:32], zll_main_word430_outR4};
  assign zll_main_word625_in = {zll_main_word626_in[97:66], zll_main_word626_in[65:0]};
  assign zll_main_word620_in = {zll_main_word625_in[97:66], zll_main_word625_in[63:32], zll_main_word625_in[31:0]};
  assign test4_in = {zll_main_word620_in[95:64], zll_main_word620_in[63:32]};
  test4  instR11 (test4_in[63:32], test4_in[31:0], extresR4[0]);
  assign zll_pure_dispatch47_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word74_in = {zll_pure_dispatch47_in[71:39], zll_pure_dispatch47_in[31:0]};
  assign zll_main_word745_in = {main_word74_in[64:32], main_word74_in[64:32], main_word74_in[31:0]};
  assign zll_main_word74_in = {zll_main_word745_in[97:65], zll_main_word745_in[31:0]};
  assign zll_main_word744_in = {zll_main_word74_in[31:0], zll_main_word74_in[64:32]};
  assign zll_main_word743_in = zll_main_word744_in[64:33];
  assign zll_main_word746_in = {zll_main_word745_in[31:0], zll_main_word745_in[64:32]};
  assign zll_main_word741_in = {zll_main_word746_in[64:33], zll_main_word746_in[31:0]};
  assign zll_main_word742_in = {zll_main_word741_in[31:0], zll_main_word741_in[63:32]};
  assign zll_pure_dispatch53_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word28_in = {zll_pure_dispatch53_in[71:39], zll_pure_dispatch53_in[31:0]};
  assign zll_main_word282_in = {main_word28_in[64:32], main_word28_in[64:32], main_word28_in[31:0]};
  assign zll_main_word283_in = {zll_main_word282_in[97:65], zll_main_word282_in[31:0]};
  assign zll_main_word28_in = {zll_main_word283_in[31:0], zll_main_word283_in[64:32]};
  assign zll_main_word281_in = zll_main_word28_in[64:33];
  assign zll_main_word286_in = {zll_main_word282_in[31:0], zll_main_word282_in[64:32]};
  assign zll_main_word284_in = {zll_main_word286_in[64:33], zll_main_word286_in[31:0]};
  assign zll_main_word285_in = {zll_main_word284_in[31:0], zll_main_word284_in[63:32]};
  assign zll_pure_dispatch31_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word38_in = {zll_pure_dispatch31_in[71:39], zll_pure_dispatch31_in[31:0]};
  assign zll_main_word385_in = {main_word38_in[64:32], main_word38_in[64:32], main_word38_in[31:0]};
  assign zll_main_word384_in = {zll_main_word385_in[97:65], zll_main_word385_in[31:0]};
  assign zll_main_word386_in = {zll_main_word384_in[31:0], zll_main_word384_in[64:32]};
  assign zll_main_word383_in = zll_main_word386_in[64:33];
  assign zll_main_word382_in = {zll_main_word385_in[31:0], zll_main_word385_in[64:32]};
  assign zll_main_word38_in = {zll_main_word382_in[64:33], zll_main_word382_in[31:0]};
  assign zll_main_word381_in = {zll_main_word38_in[31:0], zll_main_word38_in[63:32]};
  assign zll_pure_dispatch25_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word15_in = {zll_pure_dispatch25_in[71:39], zll_pure_dispatch25_in[31:0]};
  assign zll_main_word156_in = {main_word15_in[64:32], main_word15_in[64:32], main_word15_in[31:0]};
  assign zll_main_word155_in = {zll_main_word156_in[97:65], zll_main_word156_in[31:0]};
  assign zll_main_word151_in = {zll_main_word155_in[31:0], zll_main_word155_in[64:32]};
  assign zll_main_word153_in = zll_main_word151_in[64:33];
  assign zll_main_word154_in = {zll_main_word156_in[31:0], zll_main_word156_in[64:32]};
  assign zll_main_word152_in = {zll_main_word154_in[64:33], zll_main_word154_in[31:0]};
  assign zll_main_word15_in = {zll_main_word152_in[31:0], zll_main_word152_in[63:32]};
  assign zll_pure_dispatch115_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word99_in = {zll_pure_dispatch115_in[71:39], zll_pure_dispatch115_in[31:0]};
  assign zll_main_word993_in = {main_word99_in[64:32], main_word99_in[64:32], main_word99_in[31:0]};
  assign zll_main_word996_in = {zll_main_word993_in[97:65], zll_main_word993_in[31:0]};
  assign zll_main_word994_in = {zll_main_word996_in[31:0], zll_main_word996_in[64:32]};
  assign zll_main_word991_in = zll_main_word994_in[64:33];
  assign zll_main_word995_in = {zll_main_word993_in[31:0], zll_main_word993_in[64:32]};
  assign zll_main_word992_in = {zll_main_word995_in[64:33], zll_main_word995_in[31:0]};
  assign zll_main_word99_in = {zll_main_word992_in[31:0], zll_main_word992_in[63:32]};
  assign zll_pure_dispatch11_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word20_in = {zll_pure_dispatch11_in[71:39], zll_pure_dispatch11_in[31:0]};
  assign zll_main_word204_in = {main_word20_in[64:32], main_word20_in[64:32], main_word20_in[31:0]};
  assign zll_main_word202_in = {zll_main_word204_in[97:65], zll_main_word204_in[31:0]};
  assign zll_main_word201_in = {zll_main_word202_in[31:0], zll_main_word202_in[64:32]};
  assign zll_main_word205_in = zll_main_word201_in[64:33];
  assign zll_main_word20_in = {zll_main_word204_in[31:0], zll_main_word204_in[64:32]};
  assign zll_main_word203_in = {zll_main_word20_in[64:33], zll_main_word20_in[31:0]};
  assign zll_main_word206_in = {zll_main_word203_in[31:0], zll_main_word203_in[63:32]};
  assign zll_pure_dispatch101_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word9_in = {zll_pure_dispatch101_in[71:39], zll_pure_dispatch101_in[31:0]};
  assign zll_main_word9_in = {main_word9_in[64:32], main_word9_in[64:32], main_word9_in[31:0]};
  assign zll_main_word917_in = {zll_main_word9_in[97:65], zll_main_word9_in[31:0]};
  assign zll_main_word910_in = {zll_main_word917_in[31:0], zll_main_word917_in[64:32]};
  assign zll_main_word92_in = zll_main_word910_in[64:33];
  assign zll_main_word918_in = {zll_main_word9_in[31:0], zll_main_word9_in[64:32]};
  assign zll_main_word919_in = {zll_main_word918_in[64:33], zll_main_word918_in[31:0]};
  assign zll_main_word920_in = {zll_main_word919_in[31:0], zll_main_word919_in[63:32]};
  assign zll_pure_dispatch18_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word14_in = {zll_pure_dispatch18_in[71:39], zll_pure_dispatch18_in[31:0]};
  assign zll_main_word142_in = {main_word14_in[64:32], main_word14_in[64:32], main_word14_in[31:0]};
  assign zll_main_word148_in = {zll_main_word142_in[97:65], zll_main_word142_in[31:0]};
  assign zll_main_word143_in = {zll_main_word148_in[31:0], zll_main_word148_in[64:32]};
  assign zll_main_word146_in = zll_main_word143_in[64:33];
  assign zll_main_word141_in = {zll_main_word142_in[31:0], zll_main_word142_in[64:32]};
  assign zll_main_word144_in = {zll_main_word141_in[64:33], zll_main_word141_in[31:0]};
  assign zll_main_word145_in = {zll_main_word144_in[31:0], zll_main_word144_in[63:32]};
  assign zll_pure_dispatch81_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word29_in = {zll_pure_dispatch81_in[71:39], zll_pure_dispatch81_in[31:0]};
  assign zll_main_word295_in = {main_word29_in[64:32], main_word29_in[64:32], main_word29_in[31:0]};
  assign zll_main_word291_in = {zll_main_word295_in[97:65], zll_main_word295_in[31:0]};
  assign zll_main_word292_in = {zll_main_word291_in[31:0], zll_main_word291_in[64:32]};
  assign zll_main_word29_in = zll_main_word292_in[64:33];
  assign zll_main_word293_in = {zll_main_word295_in[31:0], zll_main_word295_in[64:32]};
  assign zll_main_word296_in = {zll_main_word293_in[64:33], zll_main_word293_in[31:0]};
  assign zll_main_word294_in = {zll_main_word296_in[31:0], zll_main_word296_in[63:32]};
  assign zll_pure_dispatch108_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word95_in = {zll_pure_dispatch108_in[71:39], zll_pure_dispatch108_in[31:0]};
  assign zll_main_word953_in = {main_word95_in[64:32], main_word95_in[64:32], main_word95_in[31:0]};
  assign zll_main_word955_in = {zll_main_word953_in[97:65], zll_main_word953_in[31:0]};
  assign zll_main_word954_in = {zll_main_word955_in[31:0], zll_main_word955_in[64:32]};
  assign zll_main_word95_in = zll_main_word954_in[64:33];
  assign zll_main_word952_in = {zll_main_word953_in[31:0], zll_main_word953_in[64:32]};
  assign zll_main_word956_in = {zll_main_word952_in[64:33], zll_main_word952_in[31:0]};
  assign zll_main_word951_in = {zll_main_word956_in[31:0], zll_main_word956_in[63:32]};
  assign zll_pure_dispatch46_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word77_in = {zll_pure_dispatch46_in[71:39], zll_pure_dispatch46_in[31:0]};
  assign zll_main_word776_in = {main_word77_in[64:32], main_word77_in[64:32], main_word77_in[31:0]};
  assign zll_main_word77_in = {zll_main_word776_in[97:65], zll_main_word776_in[31:0]};
  assign zll_main_word773_in = {zll_main_word77_in[31:0], zll_main_word77_in[64:32]};
  assign zll_main_word772_in = zll_main_word773_in[64:33];
  assign zll_main_word774_in = {zll_main_word776_in[31:0], zll_main_word776_in[64:32]};
  assign zll_main_word771_in = {zll_main_word774_in[64:33], zll_main_word774_in[31:0]};
  assign zll_main_word775_in = {zll_main_word771_in[31:0], zll_main_word771_in[63:32]};
  assign zll_pure_dispatch104_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word119_in = {zll_pure_dispatch104_in[71:39], zll_pure_dispatch104_in[31:0]};
  assign zll_main_word1195_in = {main_word119_in[64:32], main_word119_in[64:32], main_word119_in[31:0]};
  assign zll_main_word1196_in = {zll_main_word1195_in[97:65], zll_main_word1195_in[31:0]};
  assign zll_main_word1191_in = {zll_main_word1196_in[31:0], zll_main_word1196_in[64:32]};
  assign zll_main_word119_in = zll_main_word1191_in[64:33];
  assign zll_main_word1192_in = {zll_main_word1195_in[31:0], zll_main_word1195_in[64:32]};
  assign zll_main_word1193_in = {zll_main_word1192_in[64:33], zll_main_word1192_in[31:0]};
  assign zll_main_word1194_in = {zll_main_word1193_in[31:0], zll_main_word1193_in[63:32]};
  assign zll_pure_dispatch3_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word63_in = {zll_pure_dispatch3_in[71:39], zll_pure_dispatch3_in[31:0]};
  assign zll_main_word631_in = {main_word63_in[64:32], main_word63_in[64:32], main_word63_in[31:0]};
  assign zll_main_word634_in = {zll_main_word631_in[97:65], zll_main_word631_in[31:0]};
  assign zll_main_word633_in = {zll_main_word634_in[31:0], zll_main_word634_in[64:32]};
  assign zll_main_word635_in = zll_main_word633_in[64:33];
  assign zll_main_word63_in = {zll_main_word631_in[31:0], zll_main_word631_in[64:32]};
  assign zll_main_word636_in = {zll_main_word63_in[64:33], zll_main_word63_in[31:0]};
  assign zll_main_word632_in = {zll_main_word636_in[31:0], zll_main_word636_in[63:32]};
  assign zll_pure_dispatch38_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word65_in = {zll_pure_dispatch38_in[71:39], zll_pure_dispatch38_in[31:0]};
  assign zll_main_word654_in = {main_word65_in[64:32], main_word65_in[64:32], main_word65_in[31:0]};
  assign zll_main_word653_in = {zll_main_word654_in[97:65], zll_main_word654_in[31:0]};
  assign zll_main_word656_in = {zll_main_word653_in[31:0], zll_main_word653_in[64:32]};
  assign zll_main_word657_in = zll_main_word656_in[64:33];
  assign zll_main_word655_in = {zll_main_word654_in[31:0], zll_main_word654_in[64:32]};
  assign zll_main_word651_in = {zll_main_word655_in[64:33], zll_main_word655_in[31:0]};
  assign zll_main_word652_in = {zll_main_word651_in[31:0], zll_main_word651_in[63:32]};
  assign zll_pure_dispatch78_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word78_in = {zll_pure_dispatch78_in[71:39], zll_pure_dispatch78_in[31:0]};
  assign zll_main_word78_in = {main_word78_in[64:32], main_word78_in[64:32], main_word78_in[31:0]};
  assign zll_main_word785_in = {zll_main_word78_in[97:65], zll_main_word78_in[31:0]};
  assign zll_main_word786_in = {zll_main_word785_in[31:0], zll_main_word785_in[64:32]};
  assign zll_main_word783_in = zll_main_word786_in[64:33];
  assign zll_main_word782_in = {zll_main_word78_in[31:0], zll_main_word78_in[64:32]};
  assign zll_main_word784_in = {zll_main_word782_in[64:33], zll_main_word782_in[31:0]};
  assign zll_main_word781_in = {zll_main_word784_in[31:0], zll_main_word784_in[63:32]};
  assign zll_pure_dispatch89_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word57_in = {zll_pure_dispatch89_in[71:39], zll_pure_dispatch89_in[31:0]};
  assign zll_main_word574_in = {main_word57_in[64:32], main_word57_in[64:32], main_word57_in[31:0]};
  assign zll_main_word571_in = {zll_main_word574_in[97:65], zll_main_word574_in[31:0]};
  assign zll_main_word573_in = {zll_main_word571_in[31:0], zll_main_word571_in[64:32]};
  assign zll_main_word575_in = zll_main_word573_in[64:33];
  assign zll_main_word57_in = {zll_main_word574_in[31:0], zll_main_word574_in[64:32]};
  assign zll_main_word572_in = {zll_main_word57_in[64:33], zll_main_word57_in[31:0]};
  assign zll_main_word576_in = {zll_main_word572_in[31:0], zll_main_word572_in[63:32]};
  assign zll_pure_dispatch14_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word121_in = {zll_pure_dispatch14_in[71:39], zll_pure_dispatch14_in[31:0]};
  assign zll_main_word12111_in = {main_word121_in[64:32], main_word121_in[64:32], main_word121_in[31:0]};
  assign zll_main_word1214_in = {zll_main_word12111_in[97:65], zll_main_word12111_in[31:0]};
  assign zll_main_word1212_in = {zll_main_word1214_in[31:0], zll_main_word1214_in[64:32]};
  assign zll_main_word12110_in = zll_main_word1212_in[64:33];
  assign zll_main_word1217_in = {zll_main_word12111_in[31:0], zll_main_word12111_in[64:32]};
  assign zll_main_word1216_in = {zll_main_word1217_in[64:33], zll_main_word1217_in[31:0]};
  assign zll_main_word1218_in = {zll_main_word1216_in[31:0], zll_main_word1216_in[63:32]};
  assign zll_pure_dispatch106_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word40_in = {zll_pure_dispatch106_in[71:39], zll_pure_dispatch106_in[31:0]};
  assign zll_main_word40_in = {main_word40_in[64:32], main_word40_in[64:32], main_word40_in[31:0]};
  assign zll_main_word403_in = {zll_main_word40_in[97:65], zll_main_word40_in[31:0]};
  assign zll_main_word402_in = {zll_main_word403_in[31:0], zll_main_word403_in[64:32]};
  assign zll_main_word404_in = zll_main_word402_in[64:33];
  assign zll_main_word401_in = {zll_main_word40_in[31:0], zll_main_word40_in[64:32]};
  assign zll_main_word406_in = {zll_main_word401_in[64:33], zll_main_word401_in[31:0]};
  assign zll_main_word405_in = {zll_main_word406_in[31:0], zll_main_word406_in[63:32]};
  assign zll_pure_dispatch70_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word67_in = {zll_pure_dispatch70_in[71:39], zll_pure_dispatch70_in[31:0]};
  assign zll_main_word671_in = {main_word67_in[64:32], main_word67_in[64:32], main_word67_in[31:0]};
  assign zll_main_word673_in = {zll_main_word671_in[97:65], zll_main_word671_in[31:0]};
  assign zll_main_word676_in = {zll_main_word673_in[31:0], zll_main_word673_in[64:32]};
  assign zll_main_word67_in = zll_main_word676_in[64:33];
  assign zll_main_word674_in = {zll_main_word671_in[31:0], zll_main_word671_in[64:32]};
  assign zll_main_word675_in = {zll_main_word674_in[64:33], zll_main_word674_in[31:0]};
  assign zll_main_word672_in = {zll_main_word675_in[31:0], zll_main_word675_in[63:32]};
  assign zll_pure_dispatch39_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word33_in = {zll_pure_dispatch39_in[71:39], zll_pure_dispatch39_in[31:0]};
  assign zll_main_word335_in = {main_word33_in[64:32], main_word33_in[64:32], main_word33_in[31:0]};
  assign zll_main_word338_in = {zll_main_word335_in[97:65], zll_main_word335_in[31:0]};
  assign zll_main_word332_in = {zll_main_word338_in[31:0], zll_main_word338_in[64:32]};
  assign zll_main_word336_in = zll_main_word332_in[64:33];
  assign zll_main_word334_in = {zll_main_word335_in[31:0], zll_main_word335_in[64:32]};
  assign zll_main_word333_in = {zll_main_word334_in[64:33], zll_main_word334_in[31:0]};
  assign zll_main_word331_in = {zll_main_word333_in[31:0], zll_main_word333_in[63:32]};
  assign zll_pure_dispatch84_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word22_in = {zll_pure_dispatch84_in[71:39], zll_pure_dispatch84_in[31:0]};
  assign zll_main_word228_in = {main_word22_in[64:32], main_word22_in[64:32], main_word22_in[31:0]};
  assign zll_main_word223_in = {zll_main_word228_in[97:65], zll_main_word228_in[31:0]};
  assign zll_main_word222_in = {zll_main_word223_in[31:0], zll_main_word223_in[64:32]};
  assign zll_main_word229_in = zll_main_word222_in[64:33];
  assign zll_main_word22_in = {zll_main_word228_in[31:0], zll_main_word228_in[64:32]};
  assign zll_main_word224_in = {zll_main_word22_in[64:33], zll_main_word22_in[31:0]};
  assign zll_main_word221_in = {zll_main_word224_in[31:0], zll_main_word224_in[63:32]};
  assign zll_pure_dispatch60_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word93_in = {zll_pure_dispatch60_in[71:39], zll_pure_dispatch60_in[31:0]};
  assign zll_main_word932_in = {main_word93_in[64:32], main_word93_in[64:32], main_word93_in[31:0]};
  assign zll_main_word933_in = {zll_main_word932_in[97:65], zll_main_word932_in[31:0]};
  assign zll_main_word934_in = {zll_main_word933_in[31:0], zll_main_word933_in[64:32]};
  assign zll_main_word93_in = zll_main_word934_in[64:33];
  assign zll_main_word935_in = {zll_main_word932_in[31:0], zll_main_word932_in[64:32]};
  assign zll_main_word931_in = {zll_main_word935_in[64:33], zll_main_word935_in[31:0]};
  assign zll_main_word936_in = {zll_main_word931_in[31:0], zll_main_word931_in[63:32]};
  assign zll_pure_dispatch105_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word36_in = {zll_pure_dispatch105_in[71:39], zll_pure_dispatch105_in[31:0]};
  assign zll_main_word365_in = {main_word36_in[64:32], main_word36_in[64:32], main_word36_in[31:0]};
  assign zll_main_word362_in = {zll_main_word365_in[97:65], zll_main_word365_in[31:0]};
  assign zll_main_word361_in = {zll_main_word362_in[31:0], zll_main_word362_in[64:32]};
  assign zll_main_word366_in = zll_main_word361_in[64:33];
  assign zll_main_word36_in = {zll_main_word365_in[31:0], zll_main_word365_in[64:32]};
  assign zll_main_word363_in = {zll_main_word36_in[64:33], zll_main_word36_in[31:0]};
  assign zll_main_word364_in = {zll_main_word363_in[31:0], zll_main_word363_in[63:32]};
  assign zll_pure_dispatch107_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word110_in = {zll_pure_dispatch107_in[71:39], zll_pure_dispatch107_in[31:0]};
  assign zll_main_word1105_in = {main_word110_in[64:32], main_word110_in[64:32], main_word110_in[31:0]};
  assign zll_main_word1103_in = {zll_main_word1105_in[97:65], zll_main_word1105_in[31:0]};
  assign zll_main_word1102_in = {zll_main_word1103_in[31:0], zll_main_word1103_in[64:32]};
  assign zll_main_word1104_in = zll_main_word1102_in[64:33];
  assign zll_main_word110_in = {zll_main_word1105_in[31:0], zll_main_word1105_in[64:32]};
  assign zll_main_word1106_in = {zll_main_word110_in[64:33], zll_main_word110_in[31:0]};
  assign zll_main_word1101_in = {zll_main_word1106_in[31:0], zll_main_word1106_in[63:32]};
  assign zll_pure_dispatch109_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word84_in = {zll_pure_dispatch109_in[71:39], zll_pure_dispatch109_in[31:0]};
  assign zll_main_word841_in = {main_word84_in[64:32], main_word84_in[64:32], main_word84_in[31:0]};
  assign zll_main_word844_in = {zll_main_word841_in[97:65], zll_main_word841_in[31:0]};
  assign zll_main_word846_in = {zll_main_word844_in[31:0], zll_main_word844_in[64:32]};
  assign zll_main_word843_in = zll_main_word846_in[64:33];
  assign zll_main_word845_in = {zll_main_word841_in[31:0], zll_main_word841_in[64:32]};
  assign zll_main_word842_in = {zll_main_word845_in[64:33], zll_main_word845_in[31:0]};
  assign zll_main_word84_in = {zll_main_word842_in[31:0], zll_main_word842_in[63:32]};
  assign zll_pure_dispatch4_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word97_in = {zll_pure_dispatch4_in[71:39], zll_pure_dispatch4_in[31:0]};
  assign zll_main_word976_in = {main_word97_in[64:32], main_word97_in[64:32], main_word97_in[31:0]};
  assign zll_main_word973_in = {zll_main_word976_in[97:65], zll_main_word976_in[31:0]};
  assign zll_main_word974_in = {zll_main_word973_in[31:0], zll_main_word973_in[64:32]};
  assign zll_main_word97_in = zll_main_word974_in[64:33];
  assign zll_main_word972_in = {zll_main_word976_in[31:0], zll_main_word976_in[64:32]};
  assign zll_main_word971_in = {zll_main_word972_in[64:33], zll_main_word972_in[31:0]};
  assign zll_main_word975_in = {zll_main_word971_in[31:0], zll_main_word971_in[63:32]};
  assign zll_pure_dispatch61_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word11_in = {zll_pure_dispatch61_in[71:39], zll_pure_dispatch61_in[31:0]};
  assign zll_main_word1114_in = {main_word11_in[64:32], main_word11_in[64:32], main_word11_in[31:0]};
  assign zll_main_word1116_in = {zll_main_word1114_in[97:65], zll_main_word1114_in[31:0]};
  assign zll_main_word1117_in = {zll_main_word1116_in[31:0], zll_main_word1116_in[64:32]};
  assign zll_main_word1110_in = zll_main_word1117_in[64:33];
  assign zll_main_word1120_in = {zll_main_word1114_in[31:0], zll_main_word1114_in[64:32]};
  assign zll_main_word11_in = {zll_main_word1120_in[64:33], zll_main_word1120_in[31:0]};
  assign zll_main_word116_in = {zll_main_word11_in[31:0], zll_main_word11_in[63:32]};
  assign zll_pure_dispatch16_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word88_in = {zll_pure_dispatch16_in[71:39], zll_pure_dispatch16_in[31:0]};
  assign zll_main_word885_in = {main_word88_in[64:32], main_word88_in[64:32], main_word88_in[31:0]};
  assign zll_main_word886_in = {zll_main_word885_in[97:65], zll_main_word885_in[31:0]};
  assign zll_main_word884_in = {zll_main_word886_in[31:0], zll_main_word886_in[64:32]};
  assign zll_main_word881_in = zll_main_word884_in[64:33];
  assign zll_main_word88_in = {zll_main_word885_in[31:0], zll_main_word885_in[64:32]};
  assign zll_main_word883_in = {zll_main_word88_in[64:33], zll_main_word88_in[31:0]};
  assign zll_main_word882_in = {zll_main_word883_in[31:0], zll_main_word883_in[63:32]};
  assign zll_pure_dispatch51_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word46_in = {zll_pure_dispatch51_in[71:39], zll_pure_dispatch51_in[31:0]};
  assign zll_main_word46_in = {main_word46_in[64:32], main_word46_in[64:32], main_word46_in[31:0]};
  assign zll_main_word464_in = {zll_main_word46_in[97:65], zll_main_word46_in[31:0]};
  assign zll_main_word461_in = {zll_main_word464_in[31:0], zll_main_word464_in[64:32]};
  assign zll_main_word466_in = zll_main_word461_in[64:33];
  assign zll_main_word462_in = {zll_main_word46_in[31:0], zll_main_word46_in[64:32]};
  assign zll_main_word463_in = {zll_main_word462_in[64:33], zll_main_word462_in[31:0]};
  assign zll_main_word465_in = {zll_main_word463_in[31:0], zll_main_word463_in[63:32]};
  assign zll_pure_dispatch24_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word105_in = {zll_pure_dispatch24_in[71:39], zll_pure_dispatch24_in[31:0]};
  assign zll_main_word1054_in = {main_word105_in[64:32], main_word105_in[64:32], main_word105_in[31:0]};
  assign zll_main_word1052_in = {zll_main_word1054_in[97:65], zll_main_word1054_in[31:0]};
  assign zll_main_word1053_in = {zll_main_word1052_in[31:0], zll_main_word1052_in[64:32]};
  assign zll_main_word1051_in = zll_main_word1053_in[64:33];
  assign zll_main_word1055_in = {zll_main_word1054_in[31:0], zll_main_word1054_in[64:32]};
  assign zll_main_word105_in = {zll_main_word1055_in[64:33], zll_main_word1055_in[31:0]};
  assign zll_main_word1056_in = {zll_main_word105_in[31:0], zll_main_word105_in[63:32]};
  assign zll_pure_dispatch119_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word01_in = {zll_pure_dispatch119_in[71:39], zll_pure_dispatch119_in[31:0]};
  assign zll_main_word012_in = {main_word01_in[64:32], main_word01_in[64:32], main_word01_in[31:0]};
  assign zll_main_word011_in = {zll_main_word012_in[97:65], zll_main_word012_in[31:0]};
  assign zll_main_word010_in = {zll_main_word011_in[31:0], zll_main_word011_in[64:32]};
  assign zll_main_word08_in = zll_main_word010_in[64:33];
  assign zll_main_word01_in = {zll_main_word012_in[31:0], zll_main_word012_in[64:32]};
  assign zll_main_word07_in = {zll_main_word01_in[64:33], zll_main_word01_in[31:0]};
  assign zll_main_word04_in = {zll_main_word07_in[31:0], zll_main_word07_in[63:32]};
  assign zll_main_word06_in = zll_main_word04_in[63:32];
  ZLL_Main_word06  instR12 (zll_main_word06_in[31:0], zll_main_word06_out);
  assign zll_main_word05_in = zll_main_word06_out;
  assign zll_main_word09_inR1 = zll_main_word05_in[65:0];
  ZLL_Main_word09  instR13 (zll_main_word09_inR1[31:0], zll_main_word09_outR1);
  assign zll_pure_dispatch65_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word62_in = {zll_pure_dispatch65_in[71:39], zll_pure_dispatch65_in[31:0]};
  assign zll_main_word62_in = {main_word62_in[64:32], main_word62_in[64:32], main_word62_in[31:0]};
  assign zll_main_word627_in = {zll_main_word62_in[97:65], zll_main_word62_in[31:0]};
  assign zll_main_word621_in = {zll_main_word627_in[31:0], zll_main_word627_in[64:32]};
  assign zll_main_word628_in = zll_main_word621_in[64:33];
  assign zll_main_word624_in = {zll_main_word62_in[31:0], zll_main_word62_in[64:32]};
  assign zll_main_word623_in = {zll_main_word624_in[64:33], zll_main_word624_in[31:0]};
  assign zll_main_word622_in = {zll_main_word623_in[31:0], zll_main_word623_in[63:32]};
  assign zll_pure_dispatch55_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word2_in = {zll_pure_dispatch55_in[71:39], zll_pure_dispatch55_in[31:0]};
  assign zll_main_word226_in = {main_word2_in[64:32], main_word2_in[64:32], main_word2_in[31:0]};
  assign zll_main_word225_in = {zll_main_word226_in[97:65], zll_main_word226_in[31:0]};
  assign zll_main_word227_in = {zll_main_word225_in[31:0], zll_main_word225_in[64:32]};
  assign zll_main_word230_in = zll_main_word227_in[64:33];
  assign zll_main_word220_in = {zll_main_word226_in[31:0], zll_main_word226_in[64:32]};
  assign zll_main_word214_in = {zll_main_word220_in[64:33], zll_main_word220_in[31:0]};
  assign zll_main_word21_in = {zll_main_word214_in[31:0], zll_main_word214_in[63:32]};
  assign zll_main_word06_inR1 = zll_main_word21_in[63:32];
  ZLL_Main_word06  instR14 (zll_main_word06_inR1[31:0], zll_main_word06_outR1);
  assign zll_main_word211_in = zll_main_word06_outR1;
  assign zll_main_word314_inR1 = zll_main_word211_in[65:0];
  ZLL_Main_word314  instR15 (zll_main_word314_inR1[31:0], zll_main_word314_outR1);
  assign zll_pure_dispatch125_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word30_in = {zll_pure_dispatch125_in[71:39], zll_pure_dispatch125_in[31:0]};
  assign zll_main_word301_in = {main_word30_in[64:32], main_word30_in[64:32], main_word30_in[31:0]};
  assign zll_main_word302_in = {zll_main_word301_in[97:65], zll_main_word301_in[31:0]};
  assign zll_main_word304_in = {zll_main_word302_in[31:0], zll_main_word302_in[64:32]};
  assign zll_main_word30_in = zll_main_word304_in[64:33];
  assign zll_main_word305_in = {zll_main_word301_in[31:0], zll_main_word301_in[64:32]};
  assign zll_main_word303_in = {zll_main_word305_in[64:33], zll_main_word305_in[31:0]};
  assign zll_main_word306_in = {zll_main_word303_in[31:0], zll_main_word303_in[63:32]};
  assign zll_pure_dispatch98_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word90_in = {zll_pure_dispatch98_in[71:39], zll_pure_dispatch98_in[31:0]};
  assign zll_main_word90_in = {main_word90_in[64:32], main_word90_in[64:32], main_word90_in[31:0]};
  assign zll_main_word902_in = {zll_main_word90_in[97:65], zll_main_word90_in[31:0]};
  assign zll_main_word905_in = {zll_main_word902_in[31:0], zll_main_word902_in[64:32]};
  assign zll_main_word901_in = zll_main_word905_in[64:33];
  assign zll_main_word906_in = {zll_main_word90_in[31:0], zll_main_word90_in[64:32]};
  assign zll_main_word904_in = {zll_main_word906_in[64:33], zll_main_word906_in[31:0]};
  assign zll_main_word903_in = {zll_main_word904_in[31:0], zll_main_word904_in[63:32]};
  assign zll_pure_dispatch29_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word109_in = {zll_pure_dispatch29_in[71:39], zll_pure_dispatch29_in[31:0]};
  assign zll_main_word109_in = {main_word109_in[64:32], main_word109_in[64:32], main_word109_in[31:0]};
  assign zll_main_word1093_in = {zll_main_word109_in[97:65], zll_main_word109_in[31:0]};
  assign zll_main_word1091_in = {zll_main_word1093_in[31:0], zll_main_word1093_in[64:32]};
  assign zll_main_word1095_in = zll_main_word1091_in[64:33];
  assign zll_main_word1094_in = {zll_main_word109_in[31:0], zll_main_word109_in[64:32]};
  assign zll_main_word1096_in = {zll_main_word1094_in[64:33], zll_main_word1094_in[31:0]};
  assign zll_main_word1092_in = {zll_main_word1096_in[31:0], zll_main_word1096_in[63:32]};
  assign zll_pure_dispatch100_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word34_in = {zll_pure_dispatch100_in[71:39], zll_pure_dispatch100_in[31:0]};
  assign zll_main_word344_in = {main_word34_in[64:32], main_word34_in[64:32], main_word34_in[31:0]};
  assign zll_main_word342_in = {zll_main_word344_in[97:65], zll_main_word344_in[31:0]};
  assign zll_main_word343_in = {zll_main_word342_in[31:0], zll_main_word342_in[64:32]};
  assign zll_main_word341_in = zll_main_word343_in[64:33];
  assign zll_main_word346_in = {zll_main_word344_in[31:0], zll_main_word344_in[64:32]};
  assign zll_main_word345_in = {zll_main_word346_in[64:33], zll_main_word346_in[31:0]};
  assign zll_main_word34_in = {zll_main_word345_in[31:0], zll_main_word345_in[63:32]};
  assign zll_pure_dispatch121_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word108_in = {zll_pure_dispatch121_in[71:39], zll_pure_dispatch121_in[31:0]};
  assign zll_main_word1082_in = {main_word108_in[64:32], main_word108_in[64:32], main_word108_in[31:0]};
  assign zll_main_word1085_in = {zll_main_word1082_in[97:65], zll_main_word1082_in[31:0]};
  assign zll_main_word1086_in = {zll_main_word1085_in[31:0], zll_main_word1085_in[64:32]};
  assign zll_main_word1087_in = zll_main_word1086_in[64:33];
  assign zll_main_word1083_in = {zll_main_word1082_in[31:0], zll_main_word1082_in[64:32]};
  assign zll_main_word1081_in = {zll_main_word1083_in[64:33], zll_main_word1083_in[31:0]};
  assign zll_main_word1084_in = {zll_main_word1081_in[31:0], zll_main_word1081_in[63:32]};
  assign zll_pure_dispatch40_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word44_in = {zll_pure_dispatch40_in[71:39], zll_pure_dispatch40_in[31:0]};
  assign zll_main_word44_in = {main_word44_in[64:32], main_word44_in[64:32], main_word44_in[31:0]};
  assign zll_main_word446_in = {zll_main_word44_in[97:65], zll_main_word44_in[31:0]};
  assign zll_main_word441_in = {zll_main_word446_in[31:0], zll_main_word446_in[64:32]};
  assign zll_main_word444_in = zll_main_word441_in[64:33];
  assign zll_main_word445_in = {zll_main_word44_in[31:0], zll_main_word44_in[64:32]};
  assign zll_main_word442_in = {zll_main_word445_in[64:33], zll_main_word445_in[31:0]};
  assign zll_main_word443_in = {zll_main_word442_in[31:0], zll_main_word442_in[63:32]};
  assign zll_pure_dispatch30_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word64_in = {zll_pure_dispatch30_in[71:39], zll_pure_dispatch30_in[31:0]};
  assign zll_main_word641_in = {main_word64_in[64:32], main_word64_in[64:32], main_word64_in[31:0]};
  assign zll_main_word643_in = {zll_main_word641_in[97:65], zll_main_word641_in[31:0]};
  assign zll_main_word642_in = {zll_main_word643_in[31:0], zll_main_word643_in[64:32]};
  assign zll_main_word645_in = zll_main_word642_in[64:33];
  assign zll_main_word646_in = {zll_main_word641_in[31:0], zll_main_word641_in[64:32]};
  assign zll_main_word644_in = {zll_main_word646_in[64:33], zll_main_word646_in[31:0]};
  assign zll_main_word647_in = {zll_main_word644_in[31:0], zll_main_word644_in[63:32]};
  assign zll_pure_dispatch120_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word49_in = {zll_pure_dispatch120_in[71:39], zll_pure_dispatch120_in[31:0]};
  assign zll_main_word496_in = {main_word49_in[64:32], main_word49_in[64:32], main_word49_in[31:0]};
  assign zll_main_word491_in = {zll_main_word496_in[97:65], zll_main_word496_in[31:0]};
  assign zll_main_word495_in = {zll_main_word491_in[31:0], zll_main_word491_in[64:32]};
  assign zll_main_word494_in = zll_main_word495_in[64:33];
  assign zll_main_word49_in = {zll_main_word496_in[31:0], zll_main_word496_in[64:32]};
  assign zll_main_word492_in = {zll_main_word49_in[64:33], zll_main_word49_in[31:0]};
  assign zll_main_word493_in = {zll_main_word492_in[31:0], zll_main_word492_in[63:32]};
  assign zll_pure_dispatch73_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word73_in = {zll_pure_dispatch73_in[71:39], zll_pure_dispatch73_in[31:0]};
  assign zll_main_word73_in = {main_word73_in[64:32], main_word73_in[64:32], main_word73_in[31:0]};
  assign zll_main_word734_in = {zll_main_word73_in[97:65], zll_main_word73_in[31:0]};
  assign zll_main_word733_in = {zll_main_word734_in[31:0], zll_main_word734_in[64:32]};
  assign zll_main_word736_in = zll_main_word733_in[64:33];
  assign zll_main_word735_in = {zll_main_word73_in[31:0], zll_main_word73_in[64:32]};
  assign zll_main_word731_in = {zll_main_word735_in[64:33], zll_main_word735_in[31:0]};
  assign zll_main_word732_in = {zll_main_word731_in[31:0], zll_main_word731_in[63:32]};
  assign zll_pure_dispatch23_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word114_in = {zll_pure_dispatch23_in[71:39], zll_pure_dispatch23_in[31:0]};
  assign zll_main_word1141_in = {main_word114_in[64:32], main_word114_in[64:32], main_word114_in[31:0]};
  assign zll_main_word1144_in = {zll_main_word1141_in[97:65], zll_main_word1141_in[31:0]};
  assign zll_main_word1145_in = {zll_main_word1144_in[31:0], zll_main_word1144_in[64:32]};
  assign zll_main_word1146_in = zll_main_word1145_in[64:33];
  assign zll_main_word1143_in = {zll_main_word1141_in[31:0], zll_main_word1141_in[64:32]};
  assign zll_main_word114_in = {zll_main_word1143_in[64:33], zll_main_word1143_in[31:0]};
  assign zll_main_word1142_in = {zll_main_word114_in[31:0], zll_main_word114_in[63:32]};
  assign zll_pure_dispatch43_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word124_in = {zll_pure_dispatch43_in[71:39], zll_pure_dispatch43_in[31:0]};
  assign zll_main_word1243_in = {main_word124_in[64:32], main_word124_in[64:32], main_word124_in[31:0]};
  assign zll_main_word1247_in = {zll_main_word1243_in[97:65], zll_main_word1243_in[31:0]};
  assign zll_main_word1245_in = {zll_main_word1247_in[31:0], zll_main_word1247_in[64:32]};
  assign zll_main_word1246_in = zll_main_word1245_in[64:33];
  assign zll_main_word1244_in = {zll_main_word1243_in[31:0], zll_main_word1243_in[64:32]};
  assign zll_main_word1241_in = {zll_main_word1244_in[64:33], zll_main_word1244_in[31:0]};
  assign zll_main_word1242_in = {zll_main_word1241_in[31:0], zll_main_word1241_in[63:32]};
  assign zll_pure_dispatch95_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word48_in = {zll_pure_dispatch95_in[71:39], zll_pure_dispatch95_in[31:0]};
  assign zll_main_word485_in = {main_word48_in[64:32], main_word48_in[64:32], main_word48_in[31:0]};
  assign zll_main_word483_in = {zll_main_word485_in[97:65], zll_main_word485_in[31:0]};
  assign zll_main_word486_in = {zll_main_word483_in[31:0], zll_main_word483_in[64:32]};
  assign zll_main_word481_in = zll_main_word486_in[64:33];
  assign zll_main_word48_in = {zll_main_word485_in[31:0], zll_main_word485_in[64:32]};
  assign zll_main_word482_in = {zll_main_word48_in[64:33], zll_main_word48_in[31:0]};
  assign zll_main_word484_in = {zll_main_word482_in[31:0], zll_main_word482_in[63:32]};
  assign zll_pure_dispatch75_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word117_in = {zll_pure_dispatch75_in[71:39], zll_pure_dispatch75_in[31:0]};
  assign zll_main_word1172_in = {main_word117_in[64:32], main_word117_in[64:32], main_word117_in[31:0]};
  assign zll_main_word1175_in = {zll_main_word1172_in[97:65], zll_main_word1172_in[31:0]};
  assign zll_main_word1176_in = {zll_main_word1175_in[31:0], zll_main_word1175_in[64:32]};
  assign zll_main_word1173_in = zll_main_word1176_in[64:33];
  assign zll_main_word117_in = {zll_main_word1172_in[31:0], zll_main_word1172_in[64:32]};
  assign zll_main_word1171_in = {zll_main_word117_in[64:33], zll_main_word117_in[31:0]};
  assign zll_main_word1174_in = {zll_main_word1171_in[31:0], zll_main_word1171_in[63:32]};
  assign zll_pure_dispatch52_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word92_in = {zll_pure_dispatch52_in[71:39], zll_pure_dispatch52_in[31:0]};
  assign zll_main_word925_in = {main_word92_in[64:32], main_word92_in[64:32], main_word92_in[31:0]};
  assign zll_main_word927_in = {zll_main_word925_in[97:65], zll_main_word925_in[31:0]};
  assign zll_main_word924_in = {zll_main_word927_in[31:0], zll_main_word927_in[64:32]};
  assign zll_main_word922_in = zll_main_word924_in[64:33];
  assign zll_main_word921_in = {zll_main_word925_in[31:0], zll_main_word925_in[64:32]};
  assign zll_main_word926_in = {zll_main_word921_in[64:33], zll_main_word921_in[31:0]};
  assign zll_main_word923_in = {zll_main_word926_in[31:0], zll_main_word926_in[63:32]};
  assign zll_pure_dispatch28_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word120_in = {zll_pure_dispatch28_in[71:39], zll_pure_dispatch28_in[31:0]};
  assign zll_main_word1202_in = {main_word120_in[64:32], main_word120_in[64:32], main_word120_in[31:0]};
  assign zll_main_word1201_in = {zll_main_word1202_in[97:65], zll_main_word1202_in[31:0]};
  assign zll_main_word1204_in = {zll_main_word1201_in[31:0], zll_main_word1201_in[64:32]};
  assign zll_main_word120_in = zll_main_word1204_in[64:33];
  assign zll_main_word1205_in = {zll_main_word1202_in[31:0], zll_main_word1202_in[64:32]};
  assign zll_main_word1203_in = {zll_main_word1205_in[64:33], zll_main_word1205_in[31:0]};
  assign zll_main_word1206_in = {zll_main_word1203_in[31:0], zll_main_word1203_in[63:32]};
  assign zll_pure_dispatch59_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word104_in = {zll_pure_dispatch59_in[71:39], zll_pure_dispatch59_in[31:0]};
  assign zll_main_word104_in = {main_word104_in[64:32], main_word104_in[64:32], main_word104_in[31:0]};
  assign zll_main_word1042_in = {zll_main_word104_in[97:65], zll_main_word104_in[31:0]};
  assign zll_main_word1044_in = {zll_main_word1042_in[31:0], zll_main_word1042_in[64:32]};
  assign zll_main_word1043_in = zll_main_word1044_in[64:33];
  assign zll_main_word1045_in = {zll_main_word104_in[31:0], zll_main_word104_in[64:32]};
  assign zll_main_word1046_in = {zll_main_word1045_in[64:33], zll_main_word1045_in[31:0]};
  assign zll_main_word1041_in = {zll_main_word1046_in[31:0], zll_main_word1046_in[63:32]};
  assign zll_pure_dispatch113_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word8_in = {zll_pure_dispatch113_in[71:39], zll_pure_dispatch113_in[31:0]};
  assign zll_main_word82_in = {main_word8_in[64:32], main_word8_in[64:32], main_word8_in[31:0]};
  assign zll_main_word81_in = {zll_main_word82_in[97:65], zll_main_word82_in[31:0]};
  assign zll_main_word820_in = {zll_main_word81_in[31:0], zll_main_word81_in[64:32]};
  assign zll_main_word815_in = zll_main_word820_in[64:33];
  assign zll_main_word810_in = {zll_main_word82_in[31:0], zll_main_word82_in[64:32]};
  assign zll_main_word819_in = {zll_main_word810_in[64:33], zll_main_word810_in[31:0]};
  assign zll_main_word8_in = {zll_main_word819_in[31:0], zll_main_word819_in[63:32]};
  assign zll_pure_dispatch67_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word17_in = {zll_pure_dispatch67_in[71:39], zll_pure_dispatch67_in[31:0]};
  assign zll_main_word174_in = {main_word17_in[64:32], main_word17_in[64:32], main_word17_in[31:0]};
  assign zll_main_word175_in = {zll_main_word174_in[97:65], zll_main_word174_in[31:0]};
  assign zll_main_word176_in = {zll_main_word175_in[31:0], zll_main_word175_in[64:32]};
  assign zll_main_word173_in = zll_main_word176_in[64:33];
  assign zll_main_word17_in = {zll_main_word174_in[31:0], zll_main_word174_in[64:32]};
  assign zll_main_word172_in = {zll_main_word17_in[64:33], zll_main_word17_in[31:0]};
  assign zll_main_word171_in = {zll_main_word172_in[31:0], zll_main_word172_in[63:32]};
  assign zll_pure_dispatch36_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word50_in = {zll_pure_dispatch36_in[71:39], zll_pure_dispatch36_in[31:0]};
  assign zll_main_word506_in = {main_word50_in[64:32], main_word50_in[64:32], main_word50_in[31:0]};
  assign zll_main_word502_in = {zll_main_word506_in[97:65], zll_main_word506_in[31:0]};
  assign zll_main_word505_in = {zll_main_word502_in[31:0], zll_main_word502_in[64:32]};
  assign zll_main_word504_in = zll_main_word505_in[64:33];
  assign zll_main_word501_in = {zll_main_word506_in[31:0], zll_main_word506_in[64:32]};
  assign zll_main_word503_in = {zll_main_word501_in[64:33], zll_main_word501_in[31:0]};
  assign zll_main_word50_in = {zll_main_word503_in[31:0], zll_main_word503_in[63:32]};
  assign zll_pure_dispatch34_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word56_in = {zll_pure_dispatch34_in[71:39], zll_pure_dispatch34_in[31:0]};
  assign zll_main_word56_in = {main_word56_in[64:32], main_word56_in[64:32], main_word56_in[31:0]};
  assign zll_main_word561_in = {zll_main_word56_in[97:65], zll_main_word56_in[31:0]};
  assign zll_main_word562_in = {zll_main_word561_in[31:0], zll_main_word561_in[64:32]};
  assign zll_main_word564_in = zll_main_word562_in[64:33];
  assign zll_main_word566_in = {zll_main_word56_in[31:0], zll_main_word56_in[64:32]};
  assign zll_main_word565_in = {zll_main_word566_in[64:33], zll_main_word566_in[31:0]};
  assign zll_main_word563_in = {zll_main_word565_in[31:0], zll_main_word565_in[63:32]};
  assign zll_pure_dispatch2_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word70_in = {zll_pure_dispatch2_in[71:39], zll_pure_dispatch2_in[31:0]};
  assign zll_main_word706_in = {main_word70_in[64:32], main_word70_in[64:32], main_word70_in[31:0]};
  assign zll_main_word701_in = {zll_main_word706_in[97:65], zll_main_word706_in[31:0]};
  assign zll_main_word704_in = {zll_main_word701_in[31:0], zll_main_word701_in[64:32]};
  assign zll_main_word70_in = zll_main_word704_in[64:33];
  assign zll_main_word703_in = {zll_main_word706_in[31:0], zll_main_word706_in[64:32]};
  assign zll_main_word702_in = {zll_main_word703_in[64:33], zll_main_word703_in[31:0]};
  assign zll_main_word705_in = {zll_main_word702_in[31:0], zll_main_word702_in[63:32]};
  assign zll_pure_dispatch54_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word106_in = {zll_pure_dispatch54_in[71:39], zll_pure_dispatch54_in[31:0]};
  assign zll_main_word1061_in = {main_word106_in[64:32], main_word106_in[64:32], main_word106_in[31:0]};
  assign zll_main_word1062_in = {zll_main_word1061_in[97:65], zll_main_word1061_in[31:0]};
  assign zll_main_word1066_in = {zll_main_word1062_in[31:0], zll_main_word1062_in[64:32]};
  assign zll_main_word1064_in = zll_main_word1066_in[64:33];
  assign zll_main_word1065_in = {zll_main_word1061_in[31:0], zll_main_word1061_in[64:32]};
  assign zll_main_word106_in = {zll_main_word1065_in[64:33], zll_main_word1065_in[31:0]};
  assign zll_main_word1063_in = {zll_main_word106_in[31:0], zll_main_word106_in[63:32]};
  assign zll_pure_dispatch1_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word66_in = {zll_pure_dispatch1_in[71:39], zll_pure_dispatch1_in[31:0]};
  assign zll_main_word667_in = {main_word66_in[64:32], main_word66_in[64:32], main_word66_in[31:0]};
  assign zll_main_word661_in = {zll_main_word667_in[97:65], zll_main_word667_in[31:0]};
  assign zll_main_word663_in = {zll_main_word661_in[31:0], zll_main_word661_in[64:32]};
  assign zll_main_word665_in = zll_main_word663_in[64:33];
  assign zll_main_word664_in = {zll_main_word667_in[31:0], zll_main_word667_in[64:32]};
  assign zll_main_word662_in = {zll_main_word664_in[64:33], zll_main_word664_in[31:0]};
  assign zll_main_word666_in = {zll_main_word662_in[31:0], zll_main_word662_in[63:32]};
  assign zll_pure_dispatch35_in = {{__in0, __in1}, {__resumption_tag, __st0}};
  assign main_word23_in = {zll_pure_dispatch35_in[71:39], zll_pure_dispatch35_in[31:0]};
  assign zll_main_word235_in = {main_word23_in[64:32], main_word23_in[64:32], main_word23_in[31:0]};
  assign zll_main_word234_in = {zll_main_word235_in[97:65], zll_main_word235_in[31:0]};
  assign zll_main_word236_in = {zll_main_word234_in[31:0], zll_main_word234_in[64:32]};
  assign zll_main_word232_in = zll_main_word236_in[64:33];
  assign zll_main_word233_in = {zll_main_word235_in[31:0], zll_main_word235_in[64:32]};
  assign zll_main_word231_in = {zll_main_word233_in[64:33], zll_main_word233_in[31:0]};
  assign zll_main_word23_in = {zll_main_word231_in[31:0], zll_main_word231_in[63:32]};
  assign {__continue, __padding, __out0, __out1, __resumption_tag_next, __st0_next} = (zll_pure_dispatch35_in[38:32] == 7'h1) ? ((zll_main_word233_in[32] == 1'h0) ? {34'h20000017e, zll_main_word23_in[31:0]} : {34'h200000101, zll_main_word232_in[31:0]}) : ((zll_pure_dispatch1_in[38:32] == 7'h2) ? ((zll_main_word664_in[32] == 1'h0) ? {34'h200000127, zll_main_word666_in[31:0]} : {34'h200000102, zll_main_word665_in[31:0]}) : ((zll_pure_dispatch54_in[38:32] == 7'h3) ? ((zll_main_word1065_in[32] == 1'h0) ? {34'h200000174, zll_main_word1063_in[31:0]} : {34'h200000103, zll_main_word1064_in[31:0]}) : ((zll_pure_dispatch2_in[38:32] == 7'h4) ? ((zll_main_word703_in[32] == 1'h0) ? {34'h200000179, zll_main_word705_in[31:0]} : {34'h200000104, zll_main_word70_in[31:0]}) : ((zll_pure_dispatch34_in[38:32] == 7'h5) ? ((zll_main_word566_in[32] == 1'h0) ? {34'h20000012a, zll_main_word563_in[31:0]} : {34'h200000105, zll_main_word564_in[31:0]}) : ((zll_pure_dispatch36_in[38:32] == 7'h6) ? ((zll_main_word501_in[32] == 1'h0) ? {34'h20000017b, zll_main_word50_in[31:0]} : {34'h200000106, zll_main_word504_in[31:0]}) : ((zll_pure_dispatch67_in[38:32] == 7'h7) ? ((zll_main_word17_in[32] == 1'h0) ? {34'h200000170, zll_main_word171_in[31:0]} : {34'h200000107, zll_main_word173_in[31:0]}) : ((zll_pure_dispatch113_in[38:32] == 7'h8) ? ((zll_main_word810_in[32] == 1'h0) ? {34'h200000133, zll_main_word8_in[31:0]} : {34'h200000108, zll_main_word815_in[31:0]}) : ((zll_pure_dispatch59_in[38:32] == 7'h9) ? ((zll_main_word1045_in[32] == 1'h0) ? {34'h20000011c, zll_main_word1041_in[31:0]} : {34'h200000109, zll_main_word1043_in[31:0]}) : ((zll_pure_dispatch28_in[38:32] == 7'ha) ? ((zll_main_word1205_in[32] == 1'h0) ? {34'h200000129, zll_main_word1206_in[31:0]} : {34'h20000010a, zll_main_word120_in[31:0]}) : ((zll_pure_dispatch52_in[38:32] == 7'hb) ? ((zll_main_word921_in[32] == 1'h0) ? {34'h200000124, zll_main_word923_in[31:0]} : {34'h20000010b, zll_main_word922_in[31:0]}) : ((zll_pure_dispatch75_in[38:32] == 7'hc) ? ((zll_main_word117_in[32] == 1'h0) ? {34'h200000173, zll_main_word1174_in[31:0]} : {34'h20000010c, zll_main_word1173_in[31:0]}) : ((zll_pure_dispatch95_in[38:32] == 7'hd) ? ((zll_main_word48_in[32] == 1'h0) ? {34'h200000111, zll_main_word484_in[31:0]} : {34'h20000010d, zll_main_word481_in[31:0]}) : ((zll_pure_dispatch43_in[38:32] == 7'he) ? ((zll_main_word1244_in[32] == 1'h0) ? {34'h20000016e, zll_main_word1242_in[31:0]} : {34'h20000010e, zll_main_word1246_in[31:0]}) : ((zll_pure_dispatch23_in[38:32] == 7'hf) ? ((zll_main_word1143_in[32] == 1'h0) ? {34'h20000014f, zll_main_word1142_in[31:0]} : {34'h20000010f, zll_main_word1146_in[31:0]}) : ((zll_pure_dispatch73_in[38:32] == 7'h10) ? ((zll_main_word735_in[32] == 1'h0) ? {34'h200000139, zll_main_word732_in[31:0]} : {34'h200000110, zll_main_word736_in[31:0]}) : ((zll_pure_dispatch120_in[38:32] == 7'h11) ? ((zll_main_word49_in[32] == 1'h0) ? {34'h200000106, zll_main_word493_in[31:0]} : {34'h200000111, zll_main_word494_in[31:0]}) : ((zll_pure_dispatch30_in[38:32] == 7'h12) ? ((zll_main_word646_in[32] == 1'h0) ? {34'h20000012c, zll_main_word647_in[31:0]} : {34'h200000112, zll_main_word645_in[31:0]}) : ((zll_pure_dispatch40_in[38:32] == 7'h13) ? ((zll_main_word445_in[32] == 1'h0) ? {34'h200000143, zll_main_word443_in[31:0]} : {34'h200000113, zll_main_word444_in[31:0]}) : ((zll_pure_dispatch121_in[38:32] == 7'h14) ? ((zll_main_word1083_in[32] == 1'h0) ? {34'h200000116, zll_main_word1084_in[31:0]} : {34'h200000114, zll_main_word1087_in[31:0]}) : ((zll_pure_dispatch100_in[38:32] == 7'h15) ? ((zll_main_word346_in[32] == 1'h0) ? {34'h200000158, zll_main_word34_in[31:0]} : {34'h200000115, zll_main_word341_in[31:0]}) : ((zll_pure_dispatch29_in[38:32] == 7'h16) ? ((zll_main_word1094_in[32] == 1'h0) ? {34'h200000122, zll_main_word1092_in[31:0]} : {34'h200000116, zll_main_word1095_in[31:0]}) : ((zll_pure_dispatch98_in[38:32] == 7'h17) ? ((zll_main_word906_in[32] == 1'h0) ? {34'h200000149, zll_main_word903_in[31:0]} : {34'h200000117, zll_main_word901_in[31:0]}) : ((zll_pure_dispatch125_in[38:32] == 7'h18) ? ((zll_main_word305_in[32] == 1'h0) ? {34'h200000168, zll_main_word306_in[31:0]} : {34'h200000118, zll_main_word30_in[31:0]}) : ((zll_pure_dispatch55_in[38:32] == 7'h19) ? ((zll_main_word220_in[32] == 1'h0) ? zll_main_word314_outR1 : {34'h200000119, zll_main_word230_in[31:0]}) : ((zll_pure_dispatch65_in[38:32] == 7'h1a) ? ((zll_main_word624_in[32] == 1'h0) ? {34'h20000012d, zll_main_word622_in[31:0]} : {34'h20000011a, zll_main_word628_in[31:0]}) : ((zll_pure_dispatch119_in[38:32] == 7'h1b) ? ((zll_main_word01_in[32] == 1'h0) ? zll_main_word09_outR1 : {34'h20000011b, zll_main_word08_in[31:0]}) : ((zll_pure_dispatch24_in[38:32] == 7'h1c) ? ((zll_main_word1055_in[32] == 1'h0) ? {34'h200000103, zll_main_word1056_in[31:0]} : {34'h20000011c, zll_main_word1051_in[31:0]}) : ((zll_pure_dispatch51_in[38:32] == 7'h1d) ? ((zll_main_word462_in[32] == 1'h0) ? {34'h20000013e, zll_main_word465_in[31:0]} : {34'h20000011d, zll_main_word466_in[31:0]}) : ((zll_pure_dispatch16_in[38:32] == 7'h1e) ? ((zll_main_word88_in[32] == 1'h0) ? {34'h200000159, zll_main_word882_in[31:0]} : {34'h20000011e, zll_main_word881_in[31:0]}) : ((zll_pure_dispatch61_in[38:32] == 7'h1f) ? ((zll_main_word1120_in[32] == 1'h0) ? {34'h20000015f, zll_main_word116_in[31:0]} : {34'h20000011f, zll_main_word1110_in[31:0]}) : ((zll_pure_dispatch4_in[38:32] == 7'h20) ? ((zll_main_word972_in[32] == 1'h0) ? {34'h200000171, zll_main_word975_in[31:0]} : {34'h200000120, zll_main_word97_in[31:0]}) : ((zll_pure_dispatch109_in[38:32] == 7'h21) ? ((zll_main_word845_in[32] == 1'h0) ? {34'h20000014a, zll_main_word84_in[31:0]} : {34'h200000121, zll_main_word843_in[31:0]}) : ((zll_pure_dispatch107_in[38:32] == 7'h22) ? ((zll_main_word110_in[32] == 1'h0) ? {34'h20000017d, zll_main_word1101_in[31:0]} : {34'h200000122, zll_main_word1104_in[31:0]}) : ((zll_pure_dispatch105_in[38:32] == 7'h23) ? ((zll_main_word36_in[32] == 1'h0) ? {34'h20000016a, zll_main_word364_in[31:0]} : {34'h200000123, zll_main_word366_in[31:0]}) : ((zll_pure_dispatch60_in[38:32] == 7'h24) ? ((zll_main_word935_in[32] == 1'h0) ? {34'h200000157, zll_main_word936_in[31:0]} : {34'h200000124, zll_main_word93_in[31:0]}) : ((zll_pure_dispatch84_in[38:32] == 7'h25) ? ((zll_main_word22_in[32] == 1'h0) ? {34'h200000101, zll_main_word221_in[31:0]} : {34'h200000125, zll_main_word229_in[31:0]}) : ((zll_pure_dispatch39_in[38:32] == 7'h26) ? ((zll_main_word334_in[32] == 1'h0) ? {34'h200000115, zll_main_word331_in[31:0]} : {34'h200000126, zll_main_word336_in[31:0]}) : ((zll_pure_dispatch70_in[38:32] == 7'h27) ? ((zll_main_word674_in[32] == 1'h0) ? {34'h20000016b, zll_main_word672_in[31:0]} : {34'h200000127, zll_main_word67_in[31:0]}) : ((zll_pure_dispatch106_in[38:32] == 7'h28) ? ((zll_main_word401_in[32] == 1'h0) ? {34'h20000015c, zll_main_word405_in[31:0]} : {34'h200000128, zll_main_word404_in[31:0]}) : ((zll_pure_dispatch14_in[38:32] == 7'h29) ? ((zll_main_word1217_in[32] == 1'h0) ? {34'h200000177, zll_main_word1218_in[31:0]} : {34'h200000129, zll_main_word12110_in[31:0]}) : ((zll_pure_dispatch89_in[38:32] == 7'h2a) ? ((zll_main_word57_in[32] == 1'h0) ? {34'h200000169, zll_main_word576_in[31:0]} : {34'h20000012a, zll_main_word575_in[31:0]}) : ((zll_pure_dispatch78_in[38:32] == 7'h2b) ? ((zll_main_word782_in[32] == 1'h0) ? {34'h20000013b, zll_main_word781_in[31:0]} : {34'h20000012b, zll_main_word783_in[31:0]}) : ((zll_pure_dispatch38_in[38:32] == 7'h2c) ? ((zll_main_word655_in[32] == 1'h0) ? {34'h200000102, zll_main_word652_in[31:0]} : {34'h20000012c, zll_main_word657_in[31:0]}) : ((zll_pure_dispatch3_in[38:32] == 7'h2d) ? ((zll_main_word63_in[32] == 1'h0) ? {34'h200000112, zll_main_word632_in[31:0]} : {34'h20000012d, zll_main_word635_in[31:0]}) : ((zll_pure_dispatch104_in[38:32] == 7'h2e) ? ((zll_main_word1192_in[32] == 1'h0) ? {34'h20000010a, zll_main_word1194_in[31:0]} : {34'h20000012e, zll_main_word119_in[31:0]}) : ((zll_pure_dispatch46_in[38:32] == 7'h2f) ? ((zll_main_word774_in[32] == 1'h0) ? {34'h20000012b, zll_main_word775_in[31:0]} : {34'h20000012f, zll_main_word772_in[31:0]}) : ((zll_pure_dispatch108_in[38:32] == 7'h30) ? ((zll_main_word952_in[32] == 1'h0) ? {34'h20000015b, zll_main_word951_in[31:0]} : {34'h200000130, zll_main_word95_in[31:0]}) : ((zll_pure_dispatch81_in[38:32] == 7'h31) ? ((zll_main_word293_in[32] == 1'h0) ? {34'h200000118, zll_main_word294_in[31:0]} : {34'h200000131, zll_main_word29_in[31:0]}) : ((zll_pure_dispatch18_in[38:32] == 7'h32) ? ((zll_main_word141_in[32] == 1'h0) ? {34'h200000136, zll_main_word145_in[31:0]} : {34'h200000132, zll_main_word146_in[31:0]}) : ((zll_pure_dispatch101_in[38:32] == 7'h33) ? ((zll_main_word918_in[32] == 1'h0) ? {34'h20000017c, zll_main_word920_in[31:0]} : {34'h200000133, zll_main_word92_in[31:0]}) : ((zll_pure_dispatch11_in[38:32] == 7'h34) ? ((zll_main_word20_in[32] == 1'h0) ? {34'h200000162, zll_main_word206_in[31:0]} : {34'h200000134, zll_main_word205_in[31:0]}) : ((zll_pure_dispatch115_in[38:32] == 7'h35) ? ((zll_main_word995_in[32] == 1'h0) ? {34'h20000016f, zll_main_word99_in[31:0]} : {34'h200000135, zll_main_word991_in[31:0]}) : ((zll_pure_dispatch25_in[38:32] == 7'h36) ? ((zll_main_word154_in[32] == 1'h0) ? {34'h200000161, zll_main_word15_in[31:0]} : {34'h200000136, zll_main_word153_in[31:0]}) : ((zll_pure_dispatch31_in[38:32] == 7'h37) ? ((zll_main_word382_in[32] == 1'h0) ? {34'h200000163, zll_main_word381_in[31:0]} : {34'h200000137, zll_main_word383_in[31:0]}) : ((zll_pure_dispatch53_in[38:32] == 7'h38) ? ((zll_main_word286_in[32] == 1'h0) ? {34'h200000131, zll_main_word285_in[31:0]} : {34'h200000138, zll_main_word281_in[31:0]}) : ((zll_pure_dispatch47_in[38:32] == 7'h39) ? ((zll_main_word746_in[32] == 1'h0) ? {34'h200000147, zll_main_word742_in[31:0]} : {34'h200000139, zll_main_word743_in[31:0]}) : ((zll_pure_dispatch56_in[38:32] == 7'h3a) ? ((zll_main_word617_in[32] == 1'h0) ? {26'h2000000, extresR4, 7'h45, zll_main_word620_in[31:0]} : {34'h20000013a, zll_main_word611_in[31:0]}) : ((zll_pure_dispatch50_in[38:32] == 7'h3b) ? ((zll_main_word794_in[32] == 1'h0) ? {34'h200000164, zll_main_word792_in[31:0]} : {34'h20000013b, zll_main_word795_in[31:0]}) : ((zll_pure_dispatch33_in[38:32] == 7'h3c) ? ((zll_main_word722_in[32] == 1'h0) ? {34'h200000110, zll_main_word724_in[31:0]} : {34'h20000013c, zll_main_word723_in[31:0]}) : ((zll_pure_dispatch102_in[38:32] == 7'h3d) ? ((zll_main_word605_in[32] == 1'h0) ? {34'h200000172, zll_main_word601_in[31:0]} : {34'h20000013d, zll_main_word604_in[31:0]}) : ((zll_pure_dispatch83_in[38:32] == 7'h3e) ? ((zll_main_word476_in[32] == 1'h0) ? {34'h20000010d, zll_main_word475_in[31:0]} : {34'h20000013e, zll_main_word47_in[31:0]}) : ((zll_pure_dispatch126_in[38:32] == 7'h3f) ? ((zll_main_word1131_in[32] == 1'h0) ? {34'h20000010f, zll_main_word113_in[31:0]} : {34'h20000013f, zll_main_word1132_in[31:0]}) : ((zll_pure_dispatch118_in[38:32] == 7'h40) ? ((zll_main_word545_in[32] == 1'h0) ? {34'h200000156, zll_main_word544_in[31:0]} : {34'h200000140, zll_main_word542_in[31:0]}) : ((zll_pure_dispatch_in[38:32] == 7'h41) ? ((zll_main_word1161_in[32] == 1'h0) ? {34'h20000010c, zll_main_word1163_in[31:0]} : {34'h200000141, zll_main_word1162_in[31:0]}) : ((zll_pure_dispatch26_in[38:32] == 7'h42) ? ((zll_main_word431_in[32] == 1'h0) ? {34'h200000113, zll_main_word436_in[31:0]} : {34'h200000142, zll_main_word432_in[31:0]}) : ((zll_pure_dispatch112_in[38:32] == 7'h43) ? ((zll_main_word451_in[32] == 1'h0) ? {34'h20000011d, zll_main_word454_in[31:0]} : {34'h200000143, zll_main_word453_in[31:0]}) : ((zll_pure_dispatch63_in[38:32] == 7'h44) ? ((zll_main_word37_in[32] == 1'h0) ? {26'h2000000, extresR3, 7'h7a, zll_main_word3_in[31:0]} : zll_main_word314_out) : ((zll_pure_dispatch17_in[38:32] == 7'h45) ? ((zll_main_word710_in[32] == 1'h0) ? {34'h200000108, zll_main_word714_in[31:0]} : {34'h200000145, zll_main_word715_in[31:0]}) : ((zll_pure_dispatch66_in[38:32] == 7'h46) ? ((zll_main_word86_in[32] == 1'h0) ? {34'h20000014e, zll_main_word863_in[31:0]} : {34'h200000146, zll_main_word864_in[31:0]}) : ((zll_pure_dispatch6_in[38:32] == 7'h47) ? ((zll_main_word753_in[32] == 1'h0) ? {34'h20000014b, zll_main_word751_in[31:0]} : {34'h200000147, zll_main_word75_in[31:0]}) : ((zll_pure_dispatch13_in[38:32] == 7'h48) ? ((zll_main_word528_in[32] == 1'h0) ? {26'h2000000, extresR2, 7'h3a, zll_main_word514_in[31:0]} : {34'h200000148, zll_main_word517_in[31:0]}) : ((zll_pure_dispatch122_in[38:32] == 7'h49) ? ((zll_main_word911_in[32] == 1'h0) ? {34'h20000010b, zll_main_word916_in[31:0]} : {34'h200000149, zll_main_word915_in[31:0]}) : ((zll_pure_dispatch91_in[38:32] == 7'h4a) ? ((zll_main_word855_in[32] == 1'h0) ? {34'h200000146, zll_main_word851_in[31:0]} : {34'h20000014a, zll_main_word856_in[31:0]}) : ((zll_pure_dispatch62_in[38:32] == 7'h4b) ? ((zll_main_word764_in[32] == 1'h0) ? {34'h20000012f, zll_main_word766_in[31:0]} : {34'h20000014b, zll_main_word763_in[31:0]}) : ((zll_pure_dispatch103_in[38:32] == 7'h4c) ? ((zll_main_word195_in[32] == 1'h0) ? {34'h200000134, zll_main_word192_in[31:0]} : {34'h20000014c, zll_main_word19_in[31:0]}) : ((zll_pure_dispatch72_in[38:32] == 7'h4d) ? ((zll_main_word25_in[32] == 1'h0) ? {34'h200000155, zll_main_word255_in[31:0]} : {34'h20000014d, zll_main_word252_in[31:0]}) : ((zll_pure_dispatch21_in[38:32] == 7'h4e) ? ((zll_main_word872_in[32] == 1'h0) ? {34'h20000011e, zll_main_word876_in[31:0]} : {34'h20000014e, zll_main_word874_in[31:0]}) : ((zll_pure_dispatch69_in[38:32] == 7'h4f) ? ((zll_main_word1151_in[32] == 1'h0) ? {34'h200000141, zll_main_word1156_in[31:0]} : {34'h20000014f, zll_main_word1154_in[31:0]}) : ((zll_pure_dispatch64_in[38:32] == 7'h50) ? ((zll_main_word692_in[32] == 1'h0) ? {34'h200000104, zll_main_word694_in[31:0]} : {34'h200000150, zll_main_word693_in[31:0]}) : ((zll_pure_dispatch117_in[38:32] == 7'h51) ? ((zll_main_word13_in[32] == 1'h0) ? {34'h200000132, zll_main_word1310_in[31:0]} : {34'h200000151, zll_main_word134_in[31:0]}) : ((zll_pure_dispatch41_in[38:32] == 7'h52) ? ((zll_main_word836_in[32] == 1'h0) ? {34'h200000121, zll_main_word834_in[31:0]} : {34'h200000152, zll_main_word833_in[31:0]}) : ((zll_pure_dispatch27_in[38:32] == 7'h53) ? ((zll_main_word275_in[32] == 1'h0) ? {34'h200000138, zll_main_word276_in[31:0]} : {34'h200000153, zll_main_word273_in[31:0]}) : ((zll_pure_dispatch77_in[38:32] == 7'h54) ? ((zll_main_word1232_in[32] == 1'h0) ? {34'h20000010e, zll_main_word1234_in[31:0]} : {34'h200000154, zll_main_word1235_in[31:0]}) : ((zll_pure_dispatch48_in[38:32] == 7'h55) ? ((zll_main_word26_in[32] == 1'h0) ? {34'h200000153, zll_main_word262_in[31:0]} : {34'h200000155, zll_main_word261_in[31:0]}) : ((zll_pure_dispatch71_in[38:32] == 7'h56) ? ((zll_main_word553_in[32] == 1'h0) ? {34'h200000105, zll_main_word554_in[31:0]} : {34'h200000156, zll_main_word556_in[31:0]}) : ((zll_pure_dispatch19_in[38:32] == 7'h57) ? ((zll_main_word943_in[32] == 1'h0) ? {34'h200000130, zll_main_word941_in[31:0]} : {34'h200000157, zll_main_word946_in[31:0]}) : ((zll_pure_dispatch82_in[38:32] == 7'h58) ? ((zll_main_word352_in[32] == 1'h0) ? {34'h200000123, zll_main_word356_in[31:0]} : {34'h200000158, zll_main_word354_in[31:0]}) : ((zll_pure_dispatch44_in[38:32] == 7'h59) ? ((zll_main_word891_in[32] == 1'h0) ? {34'h200000117, zll_main_word893_in[31:0]} : {34'h200000159, zll_main_word895_in[31:0]}) : ((zll_pure_dispatch79_in[38:32] == 7'h5a) ? ((zll_main_word531_in[32] == 1'h0) ? {34'h200000140, zll_main_word534_in[31:0]} : {34'h20000015a, zll_main_word533_in[31:0]}) : ((zll_pure_dispatch32_in[38:32] == 7'h5b) ? ((zll_main_word965_in[32] == 1'h0) ? {34'h200000120, zll_main_word962_in[31:0]} : {34'h20000015b, zll_main_word963_in[31:0]}) : ((zll_pure_dispatch111_in[38:32] == 7'h5c) ? ((zll_main_word414_in[32] == 1'h0) ? {34'h20000015e, zll_main_word412_in[31:0]} : {34'h20000015c, zll_main_word416_in[31:0]}) : ((zll_pure_dispatch57_in[38:32] == 7'h5d) ? ((zll_main_word130_in[32] == 1'h0) ? {26'h2000000, extresR1, 7'h19, zll_main_word128_in[31:0]} : zll_main_word09_out) : ((zll_pure_dispatch87_in[38:32] == 7'h5e) ? ((zll_main_word42_in[32] == 1'h0) ? {34'h200000142, zll_main_word424_in[31:0]} : {34'h20000015e, zll_main_word4212_in[31:0]}) : ((zll_pure_dispatch80_in[38:32] == 7'h5f) ? ((zll_main_word127_in[32] == 1'h0) ? {34'h200000151, zll_main_word1213_in[31:0]} : {34'h20000015f, zll_main_word1210_in[31:0]}) : ((zll_pure_dispatch97_in[38:32] == 7'h60) ? ((zll_main_word1122_in[32] == 1'h0) ? {34'h20000013f, zll_main_word1125_in[31:0]} : {34'h200000160, zll_main_word1126_in[31:0]}) : ((zll_pure_dispatch88_in[38:32] == 7'h61) ? ((zll_main_word161_in[32] == 1'h0) ? {34'h200000107, zll_main_word16_in[31:0]} : {34'h200000161, zll_main_word165_in[31:0]}) : ((zll_pure_dispatch7_in[38:32] == 7'h62) ? ((zll_main_word2111_in[32] == 1'h0) ? {34'h200000125, zll_main_word2113_in[31:0]} : {34'h200000162, zll_main_word218_in[31:0]}) : ((zll_pure_dispatch90_in[38:32] == 7'h63) ? ((zll_main_word392_in[32] == 1'h0) ? {34'h200000128, zll_main_word396_in[31:0]} : {34'h200000163, zll_main_word391_in[31:0]}) : ((zll_pure_dispatch116_in[38:32] == 7'h64) ? ((zll_main_word806_in[32] == 1'h0) ? {34'h200000175, zll_main_word805_in[31:0]} : {34'h200000164, zll_main_word801_in[31:0]}) : ((zll_pure_dispatch8_in[38:32] == 7'h65) ? ((zll_main_word10110_in[32] == 1'h0) ? {34'h200000100, zll_main_word1013_in[31:0]} : {34'h200000165, zll_main_word1012_in[31:0]}) : ((zll_pure_dispatch86_in[38:32] == 7'h66) ? ((zll_main_word526_in[32] == 1'h0) ? {34'h20000015a, zll_main_word523_in[31:0]} : {34'h200000166, zll_main_word521_in[31:0]}) : ((zll_pure_dispatch15_in[38:32] == 7'h67) ? ((zll_main_word822_in[32] == 1'h0) ? {34'h200000152, zll_main_word827_in[31:0]} : {34'h200000167, zll_main_word825_in[31:0]}) : ((zll_pure_dispatch92_in[38:32] == 7'h68) ? ((zll_main_word31_in[32] == 1'h0) ? {34'h20000016c, zll_main_word3111_in[31:0]} : {34'h200000168, zll_main_word319_in[31:0]}) : ((zll_pure_dispatch58_in[38:32] == 7'h69) ? ((zll_main_word582_in[32] == 1'h0) ? {34'h20000016d, zll_main_word585_in[31:0]} : {34'h200000169, zll_main_word58_in[31:0]}) : ((zll_pure_dispatch93_in[38:32] == 7'h6a) ? ((zll_main_word374_in[32] == 1'h0) ? {34'h200000137, zll_main_word371_in[31:0]} : {34'h20000016a, zll_main_word375_in[31:0]}) : ((zll_pure_dispatch110_in[38:32] == 7'h6b) ? ((zll_main_word681_in[32] == 1'h0) ? {34'h200000150, zll_main_word686_in[31:0]} : {34'h20000016b, zll_main_word68_in[31:0]}) : ((zll_pure_dispatch99_in[38:32] == 7'h6c) ? ((zll_main_word323_in[32] == 1'h0) ? {34'h200000126, zll_main_word325_in[31:0]} : {34'h20000016c, zll_main_word322_in[31:0]}) : ((zll_pure_dispatch96_in[38:32] == 7'h6d) ? ((zll_main_word594_in[32] == 1'h0) ? {34'h20000013d, zll_main_word591_in[31:0]} : {34'h20000016d, zll_main_word593_in[31:0]}) : ((zll_pure_dispatch37_in[38:32] == 7'h6e) ? ((zll_main_word1256_in[32] == 1'h0) ? {34'h200000176, zll_main_word1253_in[31:0]} : {34'h20000016e, zll_main_word1251_in[31:0]}) : ((zll_pure_dispatch42_in[38:32] == 7'h6f) ? ((zll_main_word1003_in[32] == 1'h0) ? {34'h200000165, zll_main_word1001_in[31:0]} : {34'h20000016f, zll_main_word1006_in[31:0]}) : ((zll_pure_dispatch10_in[38:32] == 7'h70) ? ((zll_main_word186_in[32] == 1'h0) ? {34'h20000014c, zll_main_word181_in[31:0]} : {34'h200000170, zll_main_word18_in[31:0]}) : ((zll_pure_dispatch114_in[38:32] == 7'h71) ? ((zll_main_word982_in[32] == 1'h0) ? {34'h200000135, zll_main_word984_in[31:0]} : {34'h200000171, zll_main_word98_in[31:0]}) : ((zll_pure_dispatch76_in[38:32] == 7'h72) ? ((zll_main_word6112_in[32] == 1'h0) ? {34'h20000011a, zll_main_word6111_in[31:0]} : {34'h200000172, zll_main_word61_in[31:0]}) : ((zll_pure_dispatch49_in[38:32] == 7'h73) ? ((zll_main_word1181_in[32] == 1'h0) ? {34'h20000012e, zll_main_word1186_in[31:0]} : {34'h200000173, zll_main_word1183_in[31:0]}) : ((zll_pure_dispatch85_in[38:32] == 7'h74) ? ((zll_main_word1076_in[32] == 1'h0) ? {34'h200000114, zll_main_word1074_in[31:0]} : {34'h200000174, zll_main_word1071_in[31:0]}) : ((zll_pure_dispatch124_in[38:32] == 7'h75) ? ((zll_main_word811_in[32] == 1'h0) ? {34'h200000167, zll_main_word817_in[31:0]} : {34'h200000175, zll_main_word816_in[31:0]}) : ((zll_pure_dispatch12_in[38:32] == 7'h76) ? ((zll_main_word1263_in[32] == 1'h0) ? {34'h20000011b, zll_main_word1266_in[31:0]} : {34'h200000176, zll_main_word1264_in[31:0]}) : ((zll_pure_dispatch9_in[38:32] == 7'h77) ? ((zll_main_word1224_in[32] == 1'h0) ? {34'h200000154, zll_main_word122_in[31:0]} : {34'h200000177, zll_main_word1223_in[31:0]}) : ((zll_pure_dispatch123_in[38:32] == 7'h78) ? ((zll_main_word1035_in[32] == 1'h0) ? {34'h200000109, zll_main_word1032_in[31:0]} : {34'h200000178, zll_main_word1034_in[31:0]}) : ((zll_pure_dispatch68_in[38:32] == 7'h79) ? ((zll_main_word718_in[32] == 1'h0) ? {34'h20000013c, zll_main_word719_in[31:0]} : {34'h200000179, zll_main_word71_in[31:0]}) : ((zll_pure_dispatch45_in[38:32] == 7'h7a) ? ((zll_main_word423_in[32] == 1'h0) ? {26'h2000000, extres, 7'h48, zll_main_word418_in[31:0]} : {34'h20000017a, zll_main_word4_in[31:0]}) : ((zll_pure_dispatch5_in[38:32] == 7'h7b) ? ((zll_main_word5110_in[32] == 1'h0) ? {34'h200000166, zll_main_word51_in[31:0]} : {34'h20000017b, zll_main_word5111_in[31:0]}) : ((zll_pure_dispatch94_in[38:32] == 7'h7c) ? ((zll_main_word1015_in[32] == 1'h0) ? {34'h20000011f, zll_main_word1017_in[31:0]} : {34'h20000017c, zll_main_word10_in[31:0]}) : ((zll_pure_dispatch20_in[38:32] == 7'h7d) ? ((zll_main_word1118_in[32] == 1'h0) ? {34'h200000160, zll_main_word1111_in[31:0]} : {34'h20000017d, zll_main_word1119_in[31:0]}) : ((zll_pure_dispatch74_in[38:32] == 7'h7e) ? ((zll_main_word241_in[32] == 1'h0) ? {34'h20000014d, zll_main_word243_in[31:0]} : {34'h20000017e, zll_main_word244_in[31:0]}) : ((zll_main_word102_in[32] == 1'h0) ? {34'h200000178, zll_main_word1025_in[31:0]} : {34'h200000100, zll_main_word1021_in[31:0]}))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  initial {__resumption_tag, __st0} <= {7'h1b, {6'h20{1'h0}}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      {__resumption_tag, __st0} <= {7'h1b, {6'h20{1'h0}}};
    end else begin
      {__resumption_tag, __st0} <= {__resumption_tag_next, __st0_next};
    end
  end
endmodule

module ZLL_Main_word430 (input logic [63:0] arg0,
  output logic [65:0] res);
  logic [63:0] zll_main_word330_in;
  assign zll_main_word330_in = arg0;
  assign res = {2'h0, zll_main_word330_in[63:32], zll_main_word330_in[31:0]};
endmodule

module ZLL_Main_word09 (input logic [31:0] arg0,
  output logic [65:0] res);
  logic [31:0] zll_main_word013_in;
  assign zll_main_word013_in = arg0;
  assign res = {34'h20000015d, zll_main_word013_in[31:0]};
endmodule

module ZLL_Main_word06 (input logic [31:0] arg0,
  output logic [65:0] res);
  assign res = {{2'h1, {6'h20{1'h0}}}, arg0};
endmodule

module ZLL_Main_word314 (input logic [31:0] arg0,
  output logic [65:0] res);
  logic [31:0] zll_main_word318_in;
  assign zll_main_word318_in = arg0;
  assign res = {34'h200000144, zll_main_word318_in[31:0]};
endmodule