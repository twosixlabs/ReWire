module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [16:0] __in0,
  output logic [14:0] __out0);
  logic [90:0] zll_pure_dispatch2_in;
  logic [142:0] zll_pure_dispatch2_out;
  logic [90:0] zll_pure_dispatch7_in;
  logic [86:0] zll_main_reset7_in;
  logic [86:0] main_putins_in;
  logic [69:0] main_putins_out;
  logic [69:0] zll_main_loop87_in;
  logic [142:0] zll_main_loop87_out;
  logic [142:0] zll_main_reset31_in;
  logic [142:0] zll_main_reset30_in;
  logic [69:0] zll_main_reset6_in;
  logic [69:0] main_getpc_in;
  logic [75:0] main_getpc_out;
  logic [75:0] zll_main_loop101_in;
  logic [69:0] zll_main_loop101_out;
  logic [69:0] zll_main_loop87_inR1;
  logic [142:0] zll_main_loop87_outR1;
  logic [142:0] zll_main_reset24_in;
  logic [142:0] zll_main_reset23_in;
  logic [69:0] zll_main_reset3_in;
  logic [69:0] main_getout_in;
  logic [84:0] main_getout_out;
  logic [84:0] zll_main_loop94_in;
  logic [142:0] zll_main_loop94_out;
  logic [142:0] zll_main_reset19_in;
  logic [142:0] zll_main_reset18_in;
  logic [84:0] zll_main_reset2_in;
  logic [90:0] zll_pure_dispatch2_inR1;
  logic [142:0] zll_pure_dispatch2_outR1;
  logic [90:0] zll_pure_dispatch2_inR2;
  logic [142:0] zll_pure_dispatch2_outR2;
  logic [90:0] zll_pure_dispatch2_inR3;
  logic [142:0] zll_pure_dispatch2_outR3;
  logic [90:0] zll_pure_dispatch3_in;
  logic [86:0] zll_main_loop28_in;
  logic [86:0] main_putins_inR1;
  logic [69:0] main_putins_outR1;
  logic [69:0] zll_main_loop87_inR2;
  logic [142:0] zll_main_loop87_outR2;
  logic [142:0] zll_main_loop164_in;
  logic [142:0] zll_main_loop163_in;
  logic [69:0] zll_main_loop27_in;
  logic [69:0] main_incrpc_in;
  logic [69:0] main_incrpc_out;
  logic [69:0] zll_main_loop87_inR3;
  logic [142:0] zll_main_loop87_outR3;
  logic [142:0] zll_main_loop159_in;
  logic [142:0] zll_main_loop158_in;
  logic [69:0] zll_main_loop26_in;
  logic [69:0] main_getpc_inR1;
  logic [75:0] main_getpc_outR1;
  logic [75:0] zll_main_loop101_inR1;
  logic [69:0] zll_main_loop101_outR1;
  logic [69:0] zll_main_loop87_inR4;
  logic [142:0] zll_main_loop87_outR4;
  logic [142:0] zll_main_loop152_in;
  logic [142:0] zll_main_loop151_in;
  logic [69:0] zll_main_loop23_in;
  logic [69:0] main_getout_inR1;
  logic [84:0] main_getout_outR1;
  logic [84:0] zll_main_loop94_inR1;
  logic [142:0] zll_main_loop94_outR1;
  logic [142:0] zll_main_loop147_in;
  logic [142:0] zll_main_loop146_in;
  logic [84:0] zll_main_loop22_in;
  logic [90:0] zll_pure_dispatch2_inR4;
  logic [142:0] zll_pure_dispatch2_outR4;
  logic [90:0] zll_pure_dispatch1_in;
  logic [86:0] zll_main_loop16_in;
  logic [86:0] main_putins_inR2;
  logic [69:0] main_putins_outR2;
  logic [69:0] zll_main_loop87_inR5;
  logic [142:0] zll_main_loop87_outR5;
  logic [142:0] zll_main_loop132_in;
  logic [142:0] zll_main_loop131_in;
  logic [69:0] zll_main_loop15_in;
  logic [69:0] main_incrpc_inR1;
  logic [69:0] main_incrpc_outR1;
  logic [69:0] zll_main_loop87_inR6;
  logic [142:0] zll_main_loop87_outR6;
  logic [142:0] zll_main_loop127_in;
  logic [142:0] zll_main_loop126_in;
  logic [69:0] zll_main_loop14_in;
  logic [69:0] main_getpc_inR2;
  logic [75:0] main_getpc_outR2;
  logic [75:0] zll_main_loop101_inR2;
  logic [69:0] zll_main_loop101_outR2;
  logic [69:0] zll_main_loop87_inR7;
  logic [142:0] zll_main_loop87_outR7;
  logic [142:0] zll_main_loop120_in;
  logic [142:0] zll_main_loop119_in;
  logic [69:0] zll_main_loop11_in;
  logic [69:0] main_getout_inR2;
  logic [84:0] main_getout_outR2;
  logic [84:0] zll_main_loop94_inR2;
  logic [142:0] zll_main_loop94_outR2;
  logic [142:0] zll_main_loop115_in;
  logic [142:0] zll_main_loop114_in;
  logic [84:0] zll_main_loop10_in;
  logic [90:0] zll_pure_dispatch_in;
  logic [86:0] zll_main_loop9_in;
  logic [86:0] main_putins_inR3;
  logic [69:0] main_putins_outR3;
  logic [69:0] zll_main_loop87_inR8;
  logic [142:0] zll_main_loop87_outR8;
  logic [142:0] zll_main_loop110_in;
  logic [142:0] zll_main_loop109_in;
  logic [69:0] zll_main_loop8_in;
  logic [69:0] main_getdatain_in;
  logic [69:0] main_getins_in;
  logic [86:0] main_getins_out;
  logic [86:0] zll_main_getdatain2_in;
  logic [86:0] zll_main_getdatain_in;
  logic [16:0] main_datain_in;
  logic [16:0] zll_main_datain1_in;
  logic [77:0] zll_main_loop108_in;
  logic [77:0] zll_main_putreg21_in;
  logic [69:0] zll_main_putreg21_out;
  logic [69:0] zll_main_loop87_inR9;
  logic [142:0] zll_main_loop87_outR9;
  logic [142:0] zll_main_loop86_in;
  logic [142:0] zll_main_loop86_out;
  logic [0:0] __continue;
  logic [52:0] __padding;
  logic [3:0] __resumption_tag;
  logic [69:0] __st0;
  logic [3:0] __resumption_tag_next;
  logic [69:0] __st0_next;
  assign zll_pure_dispatch2_in = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch2  inst (zll_pure_dispatch2_in[90:74], zll_pure_dispatch2_in[69:0], zll_pure_dispatch2_out);
  assign zll_pure_dispatch7_in = {__in0, {__resumption_tag, __st0}};
  assign zll_main_reset7_in = {zll_pure_dispatch7_in[90:74], zll_pure_dispatch7_in[69:0]};
  assign main_putins_in = {zll_main_reset7_in[86:70], zll_main_reset7_in[69:0]};
  Main_putIns  instR1 (main_putins_in[86:70], main_putins_in[69:0], main_putins_out);
  assign zll_main_loop87_in = main_putins_out;
  ZLL_Main_loop87  instR2 (zll_main_loop87_in[69:0], zll_main_loop87_out);
  assign zll_main_reset31_in = zll_main_loop87_out;
  assign zll_main_reset30_in = zll_main_reset31_in[142:0];
  assign zll_main_reset6_in = zll_main_reset30_in[69:0];
  assign main_getpc_in = zll_main_reset6_in[69:0];
  Main_getPC  instR3 (main_getpc_in[69:0], main_getpc_out);
  assign zll_main_loop101_in = main_getpc_out;
  ZLL_Main_loop101  instR4 (zll_main_loop101_in[75:0], zll_main_loop101_out);
  assign zll_main_loop87_inR1 = zll_main_loop101_out;
  ZLL_Main_loop87  instR5 (zll_main_loop87_inR1[69:0], zll_main_loop87_outR1);
  assign zll_main_reset24_in = zll_main_loop87_outR1;
  assign zll_main_reset23_in = zll_main_reset24_in[142:0];
  assign zll_main_reset3_in = zll_main_reset23_in[69:0];
  assign main_getout_in = zll_main_reset3_in[69:0];
  Main_getOut  instR6 (main_getout_in[69:0], main_getout_out);
  assign zll_main_loop94_in = main_getout_out;
  ZLL_Main_loop94  instR7 (zll_main_loop94_in[84:0], zll_main_loop94_out);
  assign zll_main_reset19_in = zll_main_loop94_out;
  assign zll_main_reset18_in = zll_main_reset19_in[142:0];
  assign zll_main_reset2_in = {zll_main_reset18_in[84:70], zll_main_reset18_in[69:0]};
  assign zll_pure_dispatch2_inR1 = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch2  instR8 (zll_pure_dispatch2_inR1[90:74], zll_pure_dispatch2_inR1[69:0], zll_pure_dispatch2_outR1);
  assign zll_pure_dispatch2_inR2 = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch2  instR9 (zll_pure_dispatch2_inR2[90:74], zll_pure_dispatch2_inR2[69:0], zll_pure_dispatch2_outR2);
  assign zll_pure_dispatch2_inR3 = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch2  instR10 (zll_pure_dispatch2_inR3[90:74], zll_pure_dispatch2_inR3[69:0], zll_pure_dispatch2_outR3);
  assign zll_pure_dispatch3_in = {__in0, {__resumption_tag, __st0}};
  assign zll_main_loop28_in = {zll_pure_dispatch3_in[90:74], zll_pure_dispatch3_in[69:0]};
  assign main_putins_inR1 = {zll_main_loop28_in[86:70], zll_main_loop28_in[69:0]};
  Main_putIns  instR11 (main_putins_inR1[86:70], main_putins_inR1[69:0], main_putins_outR1);
  assign zll_main_loop87_inR2 = main_putins_outR1;
  ZLL_Main_loop87  instR12 (zll_main_loop87_inR2[69:0], zll_main_loop87_outR2);
  assign zll_main_loop164_in = zll_main_loop87_outR2;
  assign zll_main_loop163_in = zll_main_loop164_in[142:0];
  assign zll_main_loop27_in = zll_main_loop163_in[69:0];
  assign main_incrpc_in = zll_main_loop27_in[69:0];
  Main_incrPC  instR13 (main_incrpc_in[69:0], main_incrpc_out);
  assign zll_main_loop87_inR3 = main_incrpc_out;
  ZLL_Main_loop87  instR14 (zll_main_loop87_inR3[69:0], zll_main_loop87_outR3);
  assign zll_main_loop159_in = zll_main_loop87_outR3;
  assign zll_main_loop158_in = zll_main_loop159_in[142:0];
  assign zll_main_loop26_in = zll_main_loop158_in[69:0];
  assign main_getpc_inR1 = zll_main_loop26_in[69:0];
  Main_getPC  instR15 (main_getpc_inR1[69:0], main_getpc_outR1);
  assign zll_main_loop101_inR1 = main_getpc_outR1;
  ZLL_Main_loop101  instR16 (zll_main_loop101_inR1[75:0], zll_main_loop101_outR1);
  assign zll_main_loop87_inR4 = zll_main_loop101_outR1;
  ZLL_Main_loop87  instR17 (zll_main_loop87_inR4[69:0], zll_main_loop87_outR4);
  assign zll_main_loop152_in = zll_main_loop87_outR4;
  assign zll_main_loop151_in = zll_main_loop152_in[142:0];
  assign zll_main_loop23_in = zll_main_loop151_in[69:0];
  assign main_getout_inR1 = zll_main_loop23_in[69:0];
  Main_getOut  instR18 (main_getout_inR1[69:0], main_getout_outR1);
  assign zll_main_loop94_inR1 = main_getout_outR1;
  ZLL_Main_loop94  instR19 (zll_main_loop94_inR1[84:0], zll_main_loop94_outR1);
  assign zll_main_loop147_in = zll_main_loop94_outR1;
  assign zll_main_loop146_in = zll_main_loop147_in[142:0];
  assign zll_main_loop22_in = {zll_main_loop146_in[84:70], zll_main_loop146_in[69:0]};
  assign zll_pure_dispatch2_inR4 = {__in0, {__resumption_tag, __st0}};
  ZLL_Pure_dispatch2  instR20 (zll_pure_dispatch2_inR4[90:74], zll_pure_dispatch2_inR4[69:0], zll_pure_dispatch2_outR4);
  assign zll_pure_dispatch1_in = {__in0, {__resumption_tag, __st0}};
  assign zll_main_loop16_in = {zll_pure_dispatch1_in[90:74], zll_pure_dispatch1_in[69:0]};
  assign main_putins_inR2 = {zll_main_loop16_in[86:70], zll_main_loop16_in[69:0]};
  Main_putIns  instR21 (main_putins_inR2[86:70], main_putins_inR2[69:0], main_putins_outR2);
  assign zll_main_loop87_inR5 = main_putins_outR2;
  ZLL_Main_loop87  instR22 (zll_main_loop87_inR5[69:0], zll_main_loop87_outR5);
  assign zll_main_loop132_in = zll_main_loop87_outR5;
  assign zll_main_loop131_in = zll_main_loop132_in[142:0];
  assign zll_main_loop15_in = zll_main_loop131_in[69:0];
  assign main_incrpc_inR1 = zll_main_loop15_in[69:0];
  Main_incrPC  instR23 (main_incrpc_inR1[69:0], main_incrpc_outR1);
  assign zll_main_loop87_inR6 = main_incrpc_outR1;
  ZLL_Main_loop87  instR24 (zll_main_loop87_inR6[69:0], zll_main_loop87_outR6);
  assign zll_main_loop127_in = zll_main_loop87_outR6;
  assign zll_main_loop126_in = zll_main_loop127_in[142:0];
  assign zll_main_loop14_in = zll_main_loop126_in[69:0];
  assign main_getpc_inR2 = zll_main_loop14_in[69:0];
  Main_getPC  instR25 (main_getpc_inR2[69:0], main_getpc_outR2);
  assign zll_main_loop101_inR2 = main_getpc_outR2;
  ZLL_Main_loop101  instR26 (zll_main_loop101_inR2[75:0], zll_main_loop101_outR2);
  assign zll_main_loop87_inR7 = zll_main_loop101_outR2;
  ZLL_Main_loop87  instR27 (zll_main_loop87_inR7[69:0], zll_main_loop87_outR7);
  assign zll_main_loop120_in = zll_main_loop87_outR7;
  assign zll_main_loop119_in = zll_main_loop120_in[142:0];
  assign zll_main_loop11_in = zll_main_loop119_in[69:0];
  assign main_getout_inR2 = zll_main_loop11_in[69:0];
  Main_getOut  instR28 (main_getout_inR2[69:0], main_getout_outR2);
  assign zll_main_loop94_inR2 = main_getout_outR2;
  ZLL_Main_loop94  instR29 (zll_main_loop94_inR2[84:0], zll_main_loop94_outR2);
  assign zll_main_loop115_in = zll_main_loop94_outR2;
  assign zll_main_loop114_in = zll_main_loop115_in[142:0];
  assign zll_main_loop10_in = {zll_main_loop114_in[84:70], zll_main_loop114_in[69:0]};
  assign zll_pure_dispatch_in = {__in0, {__resumption_tag, __st0}};
  assign zll_main_loop9_in = {zll_pure_dispatch_in[90:74], zll_pure_dispatch_in[69:0]};
  assign main_putins_inR3 = {zll_main_loop9_in[86:70], zll_main_loop9_in[69:0]};
  Main_putIns  instR30 (main_putins_inR3[86:70], main_putins_inR3[69:0], main_putins_outR3);
  assign zll_main_loop87_inR8 = main_putins_outR3;
  ZLL_Main_loop87  instR31 (zll_main_loop87_inR8[69:0], zll_main_loop87_outR8);
  assign zll_main_loop110_in = zll_main_loop87_outR8;
  assign zll_main_loop109_in = zll_main_loop110_in[142:0];
  assign zll_main_loop8_in = zll_main_loop109_in[69:0];
  assign main_getdatain_in = zll_main_loop8_in[69:0];
  assign main_getins_in = main_getdatain_in[69:0];
  Main_getIns  instR32 (main_getins_in[69:0], main_getins_out);
  assign zll_main_getdatain2_in = main_getins_out;
  assign zll_main_getdatain_in = zll_main_getdatain2_in[86:0];
  assign main_datain_in = zll_main_getdatain_in[86:70];
  assign zll_main_datain1_in = main_datain_in[16:0];
  assign zll_main_loop108_in = {zll_main_datain1_in[7:0], zll_main_getdatain_in[69:0]};
  assign zll_main_putreg21_in = zll_main_loop108_in[77:0];
  ZLL_Main_putReg21  instR33 (zll_main_putreg21_in[77:70], zll_main_putreg21_in[69:0], zll_main_putreg21_out);
  assign zll_main_loop87_inR9 = zll_main_putreg21_out;
  ZLL_Main_loop87  instR34 (zll_main_loop87_inR9[69:0], zll_main_loop87_outR9);
  assign zll_main_loop86_in = zll_main_loop87_outR9;
  ZLL_Main_loop86  instR35 (zll_main_loop86_in[142:0], zll_main_loop86_out);
  assign {__continue, __padding, __out0, __resumption_tag_next, __st0_next} = (zll_pure_dispatch_in[73:70] == 4'h1) ? zll_main_loop86_out : ((zll_pure_dispatch1_in[73:70] == 4'h2) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop10_in[84:70], 4'h1, zll_main_loop10_in[69:0]} : ((zll_pure_dispatch2_inR4[73:70] == 4'h3) ? zll_pure_dispatch2_outR4 : ((zll_pure_dispatch3_in[73:70] == 4'h4) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop22_in[84:70], 4'h3, zll_main_loop22_in[69:0]} : ((zll_pure_dispatch2_inR3[73:70] == 4'h5) ? zll_pure_dispatch2_outR3 : ((zll_pure_dispatch2_inR2[73:70] == 4'h6) ? zll_pure_dispatch2_outR2 : ((zll_pure_dispatch2_inR1[73:70] == 4'h7) ? zll_pure_dispatch2_outR1 : ((zll_pure_dispatch7_in[73:70] == 4'h8) ? {{1'h1, {6'h35{1'h0}}}, zll_main_reset2_in[84:70], 4'h7, zll_main_reset2_in[69:0]} : zll_pure_dispatch2_out)))))));
  initial {__resumption_tag, __st0} <= {1'h1, {7'h49{1'h0}}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      {__resumption_tag, __st0} <= {1'h1, {7'h49{1'h0}}};
    end else begin
      {__resumption_tag, __st0} <= {__resumption_tag_next, __st0_next};
    end
  end
endmodule

module ZLL_Main_getReg5 (input logic [69:0] arg0,
  output logic [77:0] res);
  logic [139:0] zll_main_getreg10_in;
  logic [139:0] zll_main_getreg_in;
  logic [69:0] main_r0_in;
  logic [69:0] zll_main_r05_in;
  logic [61:0] zll_main_r04_in;
  logic [7:0] zll_main_r04_out;
  assign zll_main_getreg10_in = {arg0, arg0};
  assign zll_main_getreg_in = zll_main_getreg10_in[139:0];
  assign main_r0_in = zll_main_getreg_in[139:70];
  assign zll_main_r05_in = main_r0_in[69:0];
  assign zll_main_r04_in = {zll_main_r05_in[69:62], zll_main_r05_in[53:46], zll_main_r05_in[45:38], zll_main_r05_in[37:32], zll_main_r05_in[31:15], zll_main_r05_in[14:0]};
  ZLL_Main_r04  inst (zll_main_r04_in[61:54], zll_main_r04_in[53:46], zll_main_r04_in[45:38], zll_main_r04_in[37:32], zll_main_r04_in[31:15], zll_main_r04_in[14:0], zll_main_r04_out);
  assign res = {zll_main_r04_out, zll_main_getreg_in[69:0]};
endmodule

module ZLL_Main_loop86 (input logic [142:0] arg0,
  output logic [142:0] res);
  logic [142:0] zll_main_loop_in;
  logic [69:0] main_loop_in;
  logic [69:0] main_getinstr_in;
  logic [69:0] main_getins_in;
  logic [86:0] main_getins_out;
  logic [86:0] zll_main_getinstr2_in;
  logic [86:0] zll_main_getinstr_in;
  logic [16:0] main_instrin_in;
  logic [16:0] zll_main_instrin_in;
  logic [78:0] zll_main_loop264_in;
  logic [78:0] zll_main_loop262_in;
  logic [142:0] zll_main_loop261_in;
  logic [142:0] zll_main_loop260_in;
  logic [78:0] zll_main_loop61_in;
  logic [139:0] zll_main_loop259_in;
  logic [139:0] zll_main_loop257_in;
  logic [151:0] zll_main_loop256_in;
  logic [151:0] zll_main_loop254_in;
  logic [148:0] zll_main_loop53_in;
  logic [78:0] zll_main_loop217_in;
  logic [75:0] zll_main_loop216_in;
  logic [75:0] zll_main_loop60_in;
  logic [69:0] zll_main_getreg5_in;
  logic [77:0] zll_main_getreg5_out;
  logic [83:0] zll_main_loop253_in;
  logic [83:0] zll_main_loop51_in;
  logic [15:0] binop_in;
  logic [15:0] binop_inR1;
  logic [76:0] zll_main_loop84_in;
  logic [75:0] zll_main_loop83_in;
  logic [75:0] main_putpc_in;
  logic [69:0] main_putpc_out;
  logic [70:0] zll_main_loop41_in;
  logic [69:0] main_incrpc_in;
  logic [69:0] main_incrpc_out;
  logic [69:0] zll_main_loop87_in;
  logic [142:0] zll_main_loop87_out;
  logic [142:0] zll_main_loop247_in;
  logic [142:0] zll_main_loop246_in;
  logic [69:0] zll_main_loop50_in;
  logic [69:0] main_getpc_in;
  logic [75:0] main_getpc_out;
  logic [75:0] zll_main_loop101_in;
  logic [69:0] zll_main_loop101_out;
  logic [69:0] zll_main_loop87_inR1;
  logic [142:0] zll_main_loop87_outR1;
  logic [142:0] zll_main_loop201_in;
  logic [142:0] zll_main_loop200_in;
  logic [69:0] zll_main_loop47_in;
  logic [69:0] main_getout_in;
  logic [84:0] main_getout_out;
  logic [84:0] zll_main_loop94_in;
  logic [142:0] zll_main_loop94_out;
  logic [142:0] zll_main_loop196_in;
  logic [142:0] zll_main_loop195_in;
  logic [84:0] zll_main_loop46_in;
  logic [78:0] zll_main_loop214_in;
  logic [75:0] zll_main_loop213_in;
  logic [75:0] zll_main_loop212_in;
  logic [75:0] zll_main_loop58_in;
  logic [75:0] zll_main_loop57_in;
  logic [71:0] main_getreg_in;
  logic [77:0] main_getreg_out;
  logic [81:0] zll_main_loop245_in;
  logic [81:0] zll_main_loop43_in;
  logic [71:0] main_getreg_inR1;
  logic [77:0] main_getreg_outR1;
  logic [87:0] zll_main_loop79_in;
  logic [87:0] zll_main_loop42_in;
  logic [15:0] binop_inR2;
  logic [7:0] unop_in;
  logic [79:0] main_putreg_in;
  logic [79:0] zll_main_putreg44_in;
  logic [77:0] zll_main_putreg43_in;
  logic [77:0] zll_main_putreg24_in;
  logic [147:0] zll_main_putreg36_in;
  logic [147:0] zll_main_putreg12_in;
  logic [77:0] zll_main_putreg15_in;
  logic [77:0] zll_main_putreg14_in;
  logic [77:0] zll_main_putreg13_in;
  logic [79:0] zll_main_putreg42_in;
  logic [77:0] zll_main_putreg41_in;
  logic [77:0] zll_main_putreg23_in;
  logic [147:0] zll_main_putreg33_in;
  logic [147:0] zll_main_putreg7_in;
  logic [77:0] zll_main_putreg10_in;
  logic [77:0] zll_main_putreg8_in;
  logic [79:0] zll_main_putreg40_in;
  logic [77:0] zll_main_putreg39_in;
  logic [77:0] zll_main_putreg22_in;
  logic [147:0] zll_main_putreg30_in;
  logic [147:0] zll_main_putreg3_in;
  logic [77:0] zll_main_putreg5_in;
  logic [77:0] zll_main_putreg4_in;
  logic [79:0] zll_main_putreg38_in;
  logic [77:0] zll_main_putreg37_in;
  logic [77:0] zll_main_putreg21_in;
  logic [69:0] zll_main_putreg21_out;
  logic [69:0] main_incrpc_inR1;
  logic [69:0] main_incrpc_outR1;
  logic [69:0] zll_main_loop87_inR2;
  logic [142:0] zll_main_loop87_outR2;
  logic [142:0] zll_main_loop239_in;
  logic [142:0] zll_main_loop238_in;
  logic [69:0] zll_main_loop40_in;
  logic [69:0] main_getpc_inR1;
  logic [75:0] main_getpc_outR1;
  logic [75:0] zll_main_loop101_inR1;
  logic [69:0] zll_main_loop101_outR1;
  logic [69:0] zll_main_loop87_inR3;
  logic [142:0] zll_main_loop87_outR3;
  logic [142:0] zll_main_loop184_in;
  logic [142:0] zll_main_loop183_in;
  logic [69:0] zll_main_loop37_in;
  logic [69:0] main_getout_inR1;
  logic [84:0] main_getout_outR1;
  logic [84:0] zll_main_loop94_inR1;
  logic [142:0] zll_main_loop94_outR1;
  logic [142:0] zll_main_loop179_in;
  logic [142:0] zll_main_loop178_in;
  logic [84:0] zll_main_loop36_in;
  logic [78:0] zll_main_loop211_in;
  logic [75:0] zll_main_loop210_in;
  logic [75:0] zll_main_loop56_in;
  logic [69:0] zll_main_getreg5_inR1;
  logic [77:0] zll_main_getreg5_outR1;
  logic [83:0] zll_main_loop237_in;
  logic [83:0] zll_main_loop33_in;
  logic [75:0] main_putaddrout_in;
  logic [69:0] main_putaddrout_out;
  logic [77:0] zll_main_loop32_in;
  logic [77:0] main_putdataout_in;
  logic [69:0] main_getout_inR2;
  logic [84:0] main_getout_outR2;
  logic [92:0] zll_main_putdataout11_in;
  logic [92:0] zll_main_putdataout_in;
  logic [22:0] zll_main_putdataout2_in;
  logic [22:0] zll_main_putdataout1_in;
  logic [84:0] main_putout_in;
  logic [69:0] main_putout_out;
  logic [69:0] main_putweout1_in;
  logic [69:0] main_getout_inR3;
  logic [84:0] main_getout_outR3;
  logic [84:0] zll_main_putweout7_in;
  logic [84:0] zll_main_putweout2_in;
  logic [14:0] zll_main_putweout3_in;
  logic [84:0] main_putout_inR1;
  logic [69:0] main_putout_outR1;
  logic [69:0] zll_main_loop87_inR4;
  logic [142:0] zll_main_loop87_outR4;
  logic [142:0] zll_main_loop231_in;
  logic [142:0] zll_main_loop230_in;
  logic [69:0] zll_main_loop30_in;
  logic [69:0] main_getout_inR4;
  logic [84:0] main_getout_outR4;
  logic [84:0] zll_main_loop94_inR2;
  logic [142:0] zll_main_loop94_outR2;
  logic [142:0] zll_main_loop169_in;
  logic [142:0] zll_main_loop168_in;
  logic [84:0] zll_main_loop29_in;
  logic [78:0] zll_main_loop209_in;
  logic [75:0] zll_main_loop208_in;
  logic [75:0] zll_main_loop55_in;
  logic [75:0] main_putaddrout_inR1;
  logic [69:0] main_putaddrout_outR1;
  logic [69:0] main_putweout_in;
  logic [69:0] main_putweout_out;
  logic [69:0] zll_main_loop87_inR5;
  logic [142:0] zll_main_loop87_outR5;
  logic [142:0] zll_main_loop224_in;
  logic [142:0] zll_main_loop223_in;
  logic [69:0] zll_main_loop18_in;
  logic [69:0] main_getout_inR5;
  logic [84:0] main_getout_outR5;
  logic [84:0] zll_main_loop94_inR3;
  logic [142:0] zll_main_loop94_outR3;
  logic [142:0] zll_main_loop137_in;
  logic [142:0] zll_main_loop136_in;
  logic [84:0] zll_main_loop17_in;
  logic [78:0] zll_main_loop207_in;
  logic [69:0] zll_main_loop54_in;
  logic [69:0] main_incrpc_inR2;
  logic [69:0] main_incrpc_outR2;
  logic [69:0] zll_main_loop87_inR6;
  logic [142:0] zll_main_loop87_outR6;
  logic [142:0] zll_main_loop219_in;
  logic [142:0] zll_main_loop218_in;
  logic [69:0] zll_main_loop6_in;
  logic [69:0] main_getpc_inR2;
  logic [75:0] main_getpc_outR2;
  logic [75:0] zll_main_loop101_inR2;
  logic [69:0] zll_main_loop101_outR2;
  logic [69:0] zll_main_loop87_inR7;
  logic [142:0] zll_main_loop87_outR7;
  logic [142:0] zll_main_loop96_in;
  logic [142:0] zll_main_loop95_in;
  logic [69:0] zll_main_loop3_in;
  logic [69:0] main_getout_inR6;
  logic [84:0] main_getout_outR6;
  logic [84:0] zll_main_loop94_inR4;
  logic [142:0] zll_main_loop94_outR4;
  logic [142:0] zll_main_loop91_in;
  logic [142:0] zll_main_loop90_in;
  logic [84:0] zll_main_loop2_in;
  assign zll_main_loop_in = arg0;
  assign main_loop_in = zll_main_loop_in[69:0];
  assign main_getinstr_in = main_loop_in[69:0];
  assign main_getins_in = main_getinstr_in[69:0];
  Main_getIns  inst (main_getins_in[69:0], main_getins_out);
  assign zll_main_getinstr2_in = main_getins_out;
  assign zll_main_getinstr_in = zll_main_getinstr2_in[86:0];
  assign main_instrin_in = zll_main_getinstr_in[86:70];
  assign zll_main_instrin_in = main_instrin_in[16:0];
  assign zll_main_loop264_in = {zll_main_instrin_in[16:8], zll_main_getinstr_in[69:0]};
  assign zll_main_loop262_in = zll_main_loop264_in[78:0];
  assign zll_main_loop261_in = {{3'h1, {6'h3d{1'h0}}}, zll_main_loop262_in[78:70], zll_main_loop262_in[69:0]};
  assign zll_main_loop260_in = zll_main_loop261_in[142:0];
  assign zll_main_loop61_in = {zll_main_loop260_in[78:70], zll_main_loop260_in[69:0]};
  assign zll_main_loop259_in = {zll_main_loop61_in[69:0], zll_main_loop61_in[69:0]};
  assign zll_main_loop257_in = zll_main_loop259_in[139:0];
  assign zll_main_loop256_in = {zll_main_loop61_in[78:70], {3'h3, zll_main_loop257_in[139:70], zll_main_loop257_in[69:0]}};
  assign zll_main_loop254_in = {zll_main_loop256_in[151:143], zll_main_loop256_in[142:0]};
  assign zll_main_loop53_in = {zll_main_loop254_in[151:143], zll_main_loop254_in[139:70], zll_main_loop254_in[69:0]};
  assign zll_main_loop217_in = {zll_main_loop53_in[69:0], zll_main_loop53_in[148:140]};
  assign zll_main_loop216_in = {zll_main_loop217_in[78:9], zll_main_loop217_in[5:0]};
  assign zll_main_loop60_in = {zll_main_loop216_in[5:0], zll_main_loop216_in[75:6]};
  assign zll_main_getreg5_in = zll_main_loop60_in[69:0];
  ZLL_Main_getReg5  instR1 (zll_main_getreg5_in[69:0], zll_main_getreg5_out);
  assign zll_main_loop253_in = {zll_main_loop60_in[75:70], zll_main_getreg5_out};
  assign zll_main_loop51_in = {zll_main_loop253_in[83:78], zll_main_loop253_in[77:0]};
  assign binop_in = {zll_main_loop51_in[77:70], 8'h00};
  assign binop_inR1 = {zll_main_loop51_in[77:70], 8'h00};
  assign zll_main_loop84_in = {zll_main_loop51_in[69:0], zll_main_loop51_in[83:78], binop_inR1[15:8] == binop_inR1[7:0]};
  assign zll_main_loop83_in = {zll_main_loop84_in[76:7], zll_main_loop84_in[6:1]};
  assign main_putpc_in = {zll_main_loop83_in[5:0], zll_main_loop83_in[75:6]};
  Main_putPC  instR2 (main_putpc_in[75:70], main_putpc_in[69:0], main_putpc_out);
  assign zll_main_loop41_in = {zll_main_loop51_in[69:0], binop_in[15:8] == binop_in[7:0]};
  assign main_incrpc_in = zll_main_loop41_in[70:1];
  Main_incrPC  instR3 (main_incrpc_in[69:0], main_incrpc_out);
  assign zll_main_loop87_in = (zll_main_loop41_in[0] == 1'h1) ? main_incrpc_out : main_putpc_out;
  ZLL_Main_loop87  instR4 (zll_main_loop87_in[69:0], zll_main_loop87_out);
  assign zll_main_loop247_in = zll_main_loop87_out;
  assign zll_main_loop246_in = zll_main_loop247_in[142:0];
  assign zll_main_loop50_in = zll_main_loop246_in[69:0];
  assign main_getpc_in = zll_main_loop50_in[69:0];
  Main_getPC  instR5 (main_getpc_in[69:0], main_getpc_out);
  assign zll_main_loop101_in = main_getpc_out;
  ZLL_Main_loop101  instR6 (zll_main_loop101_in[75:0], zll_main_loop101_out);
  assign zll_main_loop87_inR1 = zll_main_loop101_out;
  ZLL_Main_loop87  instR7 (zll_main_loop87_inR1[69:0], zll_main_loop87_outR1);
  assign zll_main_loop201_in = zll_main_loop87_outR1;
  assign zll_main_loop200_in = zll_main_loop201_in[142:0];
  assign zll_main_loop47_in = zll_main_loop200_in[69:0];
  assign main_getout_in = zll_main_loop47_in[69:0];
  Main_getOut  instR8 (main_getout_in[69:0], main_getout_out);
  assign zll_main_loop94_in = main_getout_out;
  ZLL_Main_loop94  instR9 (zll_main_loop94_in[84:0], zll_main_loop94_out);
  assign zll_main_loop196_in = zll_main_loop94_out;
  assign zll_main_loop195_in = zll_main_loop196_in[142:0];
  assign zll_main_loop46_in = {zll_main_loop195_in[84:70], zll_main_loop195_in[69:0]};
  assign zll_main_loop214_in = {zll_main_loop53_in[69:0], zll_main_loop53_in[148:140]};
  assign zll_main_loop213_in = {zll_main_loop214_in[78:9], zll_main_loop214_in[5:4], zll_main_loop214_in[3:2], zll_main_loop214_in[1:0]};
  assign zll_main_loop212_in = {zll_main_loop213_in[75:6], zll_main_loop213_in[3:2], zll_main_loop213_in[5:4], zll_main_loop213_in[1:0]};
  assign zll_main_loop58_in = {zll_main_loop212_in[3:2], zll_main_loop212_in[5:4], zll_main_loop212_in[1:0], zll_main_loop212_in[75:6]};
  assign zll_main_loop57_in = {zll_main_loop58_in[73:72], zll_main_loop58_in[75:74], zll_main_loop58_in[71:70], zll_main_loop58_in[69:0]};
  assign main_getreg_in = {zll_main_loop57_in[75:74], zll_main_loop57_in[69:0]};
  Main_getReg  instR10 (main_getreg_in[71:70], main_getreg_in[69:0], main_getreg_out);
  assign zll_main_loop245_in = {zll_main_loop57_in[71:70], zll_main_loop57_in[73:72], main_getreg_out};
  assign zll_main_loop43_in = {zll_main_loop245_in[81:80], zll_main_loop245_in[79:78], zll_main_loop245_in[77:0]};
  assign main_getreg_inR1 = {zll_main_loop43_in[81:80], zll_main_loop43_in[69:0]};
  Main_getReg  instR11 (main_getreg_inR1[71:70], main_getreg_inR1[69:0], main_getreg_outR1);
  assign zll_main_loop79_in = {zll_main_loop43_in[77:70], zll_main_loop43_in[79:78], main_getreg_outR1};
  assign zll_main_loop42_in = {zll_main_loop79_in[87:80], zll_main_loop79_in[79:78], zll_main_loop79_in[77:0]};
  assign binop_inR2 = {zll_main_loop42_in[87:80], zll_main_loop42_in[77:70]};
  assign unop_in = binop_inR2[15:8] & binop_inR2[7:0];
  assign main_putreg_in = {zll_main_loop42_in[79:78], ~unop_in[7:0], zll_main_loop42_in[69:0]};
  assign zll_main_putreg44_in = {main_putreg_in[69:0], main_putreg_in[79:78], main_putreg_in[77:70]};
  assign zll_main_putreg43_in = {zll_main_putreg44_in[79:10], zll_main_putreg44_in[7:0]};
  assign zll_main_putreg24_in = {zll_main_putreg43_in[7:0], zll_main_putreg43_in[77:8]};
  assign zll_main_putreg36_in = {zll_main_putreg24_in[77:70], zll_main_putreg24_in[69:0], zll_main_putreg24_in[69:0]};
  assign zll_main_putreg12_in = {zll_main_putreg36_in[147:140], zll_main_putreg36_in[139:0]};
  assign zll_main_putreg15_in = {zll_main_putreg12_in[147:140], zll_main_putreg12_in[139:70]};
  assign zll_main_putreg14_in = {zll_main_putreg15_in[77:70], zll_main_putreg15_in[61:54], zll_main_putreg15_in[69:62], zll_main_putreg15_in[53:46], zll_main_putreg15_in[45:38], zll_main_putreg15_in[37:32], zll_main_putreg15_in[31:15], zll_main_putreg15_in[14:0]};
  assign zll_main_putreg13_in = {zll_main_putreg14_in[77:70], zll_main_putreg14_in[69:62], zll_main_putreg14_in[53:46], zll_main_putreg14_in[61:54], zll_main_putreg14_in[45:38], zll_main_putreg14_in[37:32], zll_main_putreg14_in[31:15], zll_main_putreg14_in[14:0]};
  assign zll_main_putreg42_in = {main_putreg_in[69:0], main_putreg_in[79:78], main_putreg_in[77:70]};
  assign zll_main_putreg41_in = {zll_main_putreg42_in[79:10], zll_main_putreg42_in[7:0]};
  assign zll_main_putreg23_in = {zll_main_putreg41_in[7:0], zll_main_putreg41_in[77:8]};
  assign zll_main_putreg33_in = {zll_main_putreg23_in[77:70], zll_main_putreg23_in[69:0], zll_main_putreg23_in[69:0]};
  assign zll_main_putreg7_in = {zll_main_putreg33_in[147:140], zll_main_putreg33_in[139:0]};
  assign zll_main_putreg10_in = {zll_main_putreg7_in[147:140], zll_main_putreg7_in[139:70]};
  assign zll_main_putreg8_in = {zll_main_putreg10_in[69:62], zll_main_putreg10_in[77:70], zll_main_putreg10_in[61:54], zll_main_putreg10_in[53:46], zll_main_putreg10_in[45:38], zll_main_putreg10_in[37:32], zll_main_putreg10_in[31:15], zll_main_putreg10_in[14:0]};
  assign zll_main_putreg40_in = {main_putreg_in[69:0], main_putreg_in[79:78], main_putreg_in[77:70]};
  assign zll_main_putreg39_in = {zll_main_putreg40_in[79:10], zll_main_putreg40_in[7:0]};
  assign zll_main_putreg22_in = {zll_main_putreg39_in[7:0], zll_main_putreg39_in[77:8]};
  assign zll_main_putreg30_in = {zll_main_putreg22_in[77:70], zll_main_putreg22_in[69:0], zll_main_putreg22_in[69:0]};
  assign zll_main_putreg3_in = {zll_main_putreg30_in[147:140], zll_main_putreg30_in[139:0]};
  assign zll_main_putreg5_in = {zll_main_putreg3_in[147:140], zll_main_putreg3_in[139:70]};
  assign zll_main_putreg4_in = {zll_main_putreg5_in[69:62], zll_main_putreg5_in[77:70], zll_main_putreg5_in[61:54], zll_main_putreg5_in[53:46], zll_main_putreg5_in[45:38], zll_main_putreg5_in[37:32], zll_main_putreg5_in[31:15], zll_main_putreg5_in[14:0]};
  assign zll_main_putreg38_in = {main_putreg_in[69:0], main_putreg_in[79:78], main_putreg_in[77:70]};
  assign zll_main_putreg37_in = {zll_main_putreg38_in[79:10], zll_main_putreg38_in[7:0]};
  assign zll_main_putreg21_in = {zll_main_putreg37_in[7:0], zll_main_putreg37_in[77:8]};
  ZLL_Main_putReg21  instR12 (zll_main_putreg21_in[77:70], zll_main_putreg21_in[69:0], zll_main_putreg21_out);
  assign main_incrpc_inR1 = (zll_main_putreg38_in[9:8] == 2'h0) ? zll_main_putreg21_out : ((zll_main_putreg40_in[9:8] == 2'h1) ? {zll_main_putreg4_in[77:70], zll_main_putreg4_in[69:62], zll_main_putreg4_in[53:46], zll_main_putreg4_in[45:38], zll_main_putreg4_in[37:32], zll_main_putreg4_in[31:15], zll_main_putreg4_in[14:0]} : ((zll_main_putreg42_in[9:8] == 2'h2) ? {zll_main_putreg8_in[77:70], zll_main_putreg8_in[61:54], zll_main_putreg8_in[69:62], zll_main_putreg8_in[45:38], zll_main_putreg8_in[37:32], zll_main_putreg8_in[31:15], zll_main_putreg8_in[14:0]} : {zll_main_putreg13_in[53:46], zll_main_putreg13_in[69:62], zll_main_putreg13_in[61:54], zll_main_putreg13_in[77:70], zll_main_putreg13_in[37:32], zll_main_putreg13_in[31:15], zll_main_putreg13_in[14:0]}));
  Main_incrPC  instR13 (main_incrpc_inR1[69:0], main_incrpc_outR1);
  assign zll_main_loop87_inR2 = main_incrpc_outR1;
  ZLL_Main_loop87  instR14 (zll_main_loop87_inR2[69:0], zll_main_loop87_outR2);
  assign zll_main_loop239_in = zll_main_loop87_outR2;
  assign zll_main_loop238_in = zll_main_loop239_in[142:0];
  assign zll_main_loop40_in = zll_main_loop238_in[69:0];
  assign main_getpc_inR1 = zll_main_loop40_in[69:0];
  Main_getPC  instR15 (main_getpc_inR1[69:0], main_getpc_outR1);
  assign zll_main_loop101_inR1 = main_getpc_outR1;
  ZLL_Main_loop101  instR16 (zll_main_loop101_inR1[75:0], zll_main_loop101_outR1);
  assign zll_main_loop87_inR3 = zll_main_loop101_outR1;
  ZLL_Main_loop87  instR17 (zll_main_loop87_inR3[69:0], zll_main_loop87_outR3);
  assign zll_main_loop184_in = zll_main_loop87_outR3;
  assign zll_main_loop183_in = zll_main_loop184_in[142:0];
  assign zll_main_loop37_in = zll_main_loop183_in[69:0];
  assign main_getout_inR1 = zll_main_loop37_in[69:0];
  Main_getOut  instR18 (main_getout_inR1[69:0], main_getout_outR1);
  assign zll_main_loop94_inR1 = main_getout_outR1;
  ZLL_Main_loop94  instR19 (zll_main_loop94_inR1[84:0], zll_main_loop94_outR1);
  assign zll_main_loop179_in = zll_main_loop94_outR1;
  assign zll_main_loop178_in = zll_main_loop179_in[142:0];
  assign zll_main_loop36_in = {zll_main_loop178_in[84:70], zll_main_loop178_in[69:0]};
  assign zll_main_loop211_in = {zll_main_loop53_in[69:0], zll_main_loop53_in[148:140]};
  assign zll_main_loop210_in = {zll_main_loop211_in[78:9], zll_main_loop211_in[5:0]};
  assign zll_main_loop56_in = {zll_main_loop210_in[5:0], zll_main_loop210_in[75:6]};
  assign zll_main_getreg5_inR1 = zll_main_loop56_in[69:0];
  ZLL_Main_getReg5  instR20 (zll_main_getreg5_inR1[69:0], zll_main_getreg5_outR1);
  assign zll_main_loop237_in = {zll_main_loop56_in[75:70], zll_main_getreg5_outR1};
  assign zll_main_loop33_in = {zll_main_loop237_in[83:78], zll_main_loop237_in[77:0]};
  assign main_putaddrout_in = {zll_main_loop33_in[83:78], zll_main_loop33_in[69:0]};
  Main_putAddrOut  instR21 (main_putaddrout_in[75:70], main_putaddrout_in[69:0], main_putaddrout_out);
  assign zll_main_loop32_in = {zll_main_loop33_in[77:70], main_putaddrout_out};
  assign main_putdataout_in = {zll_main_loop32_in[77:70], zll_main_loop32_in[69:0]};
  assign main_getout_inR2 = main_putdataout_in[69:0];
  Main_getOut  instR22 (main_getout_inR2[69:0], main_getout_outR2);
  assign zll_main_putdataout11_in = {main_putdataout_in[77:70], main_getout_outR2};
  assign zll_main_putdataout_in = {zll_main_putdataout11_in[92:85], zll_main_putdataout11_in[84:0]};
  assign zll_main_putdataout2_in = {zll_main_putdataout_in[92:85], zll_main_putdataout_in[84:70]};
  assign zll_main_putdataout1_in = {zll_main_putdataout2_in[13:8], zll_main_putdataout2_in[22:15], zll_main_putdataout2_in[14], zll_main_putdataout2_in[7:0]};
  assign main_putout_in = {{zll_main_putdataout1_in[8], zll_main_putdataout1_in[22:17], zll_main_putdataout1_in[16:9]}, zll_main_putdataout_in[69:0]};
  Main_putOut  instR23 (main_putout_in[84:70], main_putout_in[69:0], main_putout_out);
  assign main_putweout1_in = main_putout_out;
  assign main_getout_inR3 = main_putweout1_in[69:0];
  Main_getOut  instR24 (main_getout_inR3[69:0], main_getout_outR3);
  assign zll_main_putweout7_in = main_getout_outR3;
  assign zll_main_putweout2_in = zll_main_putweout7_in[84:0];
  assign zll_main_putweout3_in = zll_main_putweout2_in[84:70];
  assign main_putout_inR1 = {{1'h1, zll_main_putweout3_in[13:8], zll_main_putweout3_in[7:0]}, zll_main_putweout2_in[69:0]};
  Main_putOut  instR25 (main_putout_inR1[84:70], main_putout_inR1[69:0], main_putout_outR1);
  assign zll_main_loop87_inR4 = main_putout_outR1;
  ZLL_Main_loop87  instR26 (zll_main_loop87_inR4[69:0], zll_main_loop87_outR4);
  assign zll_main_loop231_in = zll_main_loop87_outR4;
  assign zll_main_loop230_in = zll_main_loop231_in[142:0];
  assign zll_main_loop30_in = zll_main_loop230_in[69:0];
  assign main_getout_inR4 = zll_main_loop30_in[69:0];
  Main_getOut  instR27 (main_getout_inR4[69:0], main_getout_outR4);
  assign zll_main_loop94_inR2 = main_getout_outR4;
  ZLL_Main_loop94  instR28 (zll_main_loop94_inR2[84:0], zll_main_loop94_outR2);
  assign zll_main_loop169_in = zll_main_loop94_outR2;
  assign zll_main_loop168_in = zll_main_loop169_in[142:0];
  assign zll_main_loop29_in = {zll_main_loop168_in[84:70], zll_main_loop168_in[69:0]};
  assign zll_main_loop209_in = {zll_main_loop53_in[69:0], zll_main_loop53_in[148:140]};
  assign zll_main_loop208_in = {zll_main_loop209_in[78:9], zll_main_loop209_in[5:0]};
  assign zll_main_loop55_in = {zll_main_loop208_in[5:0], zll_main_loop208_in[75:6]};
  assign main_putaddrout_inR1 = {zll_main_loop55_in[75:70], zll_main_loop55_in[69:0]};
  Main_putAddrOut  instR29 (main_putaddrout_inR1[75:70], main_putaddrout_inR1[69:0], main_putaddrout_outR1);
  assign main_putweout_in = main_putaddrout_outR1;
  Main_putWeOut  instR30 (main_putweout_in[69:0], main_putweout_out);
  assign zll_main_loop87_inR5 = main_putweout_out;
  ZLL_Main_loop87  instR31 (zll_main_loop87_inR5[69:0], zll_main_loop87_outR5);
  assign zll_main_loop224_in = zll_main_loop87_outR5;
  assign zll_main_loop223_in = zll_main_loop224_in[142:0];
  assign zll_main_loop18_in = zll_main_loop223_in[69:0];
  assign main_getout_inR5 = zll_main_loop18_in[69:0];
  Main_getOut  instR32 (main_getout_inR5[69:0], main_getout_outR5);
  assign zll_main_loop94_inR3 = main_getout_outR5;
  ZLL_Main_loop94  instR33 (zll_main_loop94_inR3[84:0], zll_main_loop94_outR3);
  assign zll_main_loop137_in = zll_main_loop94_outR3;
  assign zll_main_loop136_in = zll_main_loop137_in[142:0];
  assign zll_main_loop17_in = {zll_main_loop136_in[84:70], zll_main_loop136_in[69:0]};
  assign zll_main_loop207_in = {zll_main_loop53_in[69:0], zll_main_loop53_in[148:140]};
  assign zll_main_loop54_in = zll_main_loop207_in[78:9];
  assign main_incrpc_inR2 = zll_main_loop54_in[69:0];
  Main_incrPC  instR34 (main_incrpc_inR2[69:0], main_incrpc_outR2);
  assign zll_main_loop87_inR6 = main_incrpc_outR2;
  ZLL_Main_loop87  instR35 (zll_main_loop87_inR6[69:0], zll_main_loop87_outR6);
  assign zll_main_loop219_in = zll_main_loop87_outR6;
  assign zll_main_loop218_in = zll_main_loop219_in[142:0];
  assign zll_main_loop6_in = zll_main_loop218_in[69:0];
  assign main_getpc_inR2 = zll_main_loop6_in[69:0];
  Main_getPC  instR36 (main_getpc_inR2[69:0], main_getpc_outR2);
  assign zll_main_loop101_inR2 = main_getpc_outR2;
  ZLL_Main_loop101  instR37 (zll_main_loop101_inR2[75:0], zll_main_loop101_outR2);
  assign zll_main_loop87_inR7 = zll_main_loop101_outR2;
  ZLL_Main_loop87  instR38 (zll_main_loop87_inR7[69:0], zll_main_loop87_outR7);
  assign zll_main_loop96_in = zll_main_loop87_outR7;
  assign zll_main_loop95_in = zll_main_loop96_in[142:0];
  assign zll_main_loop3_in = zll_main_loop95_in[69:0];
  assign main_getout_inR6 = zll_main_loop3_in[69:0];
  Main_getOut  instR39 (main_getout_inR6[69:0], main_getout_outR6);
  assign zll_main_loop94_inR4 = main_getout_outR6;
  ZLL_Main_loop94  instR40 (zll_main_loop94_inR4[84:0], zll_main_loop94_outR4);
  assign zll_main_loop91_in = zll_main_loop94_outR4;
  assign zll_main_loop90_in = zll_main_loop91_in[142:0];
  assign zll_main_loop2_in = {zll_main_loop90_in[84:70], zll_main_loop90_in[69:0]};
  assign res = (zll_main_loop207_in[8:6] == 3'h0) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop2_in[84:70], 4'h0, zll_main_loop2_in[69:0]} : ((zll_main_loop209_in[8:6] == 3'h1) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop17_in[84:70], 4'h2, zll_main_loop17_in[69:0]} : ((zll_main_loop211_in[8:6] == 3'h2) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop29_in[84:70], 4'h4, zll_main_loop29_in[69:0]} : ((zll_main_loop214_in[8:6] == 3'h3) ? {{1'h1, {6'h35{1'h0}}}, zll_main_loop36_in[84:70], 4'h5, zll_main_loop36_in[69:0]} : {{1'h1, {6'h35{1'h0}}}, zll_main_loop46_in[84:70], 4'h6, zll_main_loop46_in[69:0]})));
endmodule

module ZLL_Main_loop87 (input logic [69:0] arg0,
  output logic [142:0] res);
  assign res = {{7'h49{1'h0}}, arg0};
endmodule

module ZLL_Main_loop94 (input logic [84:0] arg0,
  output logic [142:0] res);
  logic [84:0] zll_main_loop92_in;
  assign zll_main_loop92_in = arg0;
  assign res = {{2'h1, {6'h38{1'h0}}}, zll_main_loop92_in[84:70], zll_main_loop92_in[69:0]};
endmodule

module ZLL_Main_loop101 (input logic [75:0] arg0,
  output logic [69:0] res);
  logic [75:0] zll_main_loop5_in;
  logic [75:0] main_putaddrout_in;
  logic [69:0] main_putaddrout_out;
  logic [69:0] main_putweout_in;
  logic [69:0] main_putweout_out;
  assign zll_main_loop5_in = arg0;
  assign main_putaddrout_in = {zll_main_loop5_in[75:70], zll_main_loop5_in[69:0]};
  Main_putAddrOut  inst (main_putaddrout_in[75:70], main_putaddrout_in[69:0], main_putaddrout_out);
  assign main_putweout_in = main_putaddrout_out;
  Main_putWeOut  instR1 (main_putweout_in[69:0], main_putweout_out);
  assign res = main_putweout_out;
endmodule

module ZLL_Main_putReg21 (input logic [7:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [147:0] zll_main_putreg27_in;
  logic [147:0] zll_main_putreg_in;
  logic [77:0] zll_main_putreg1_in;
  assign zll_main_putreg27_in = {arg0, arg1, arg1};
  assign zll_main_putreg_in = {zll_main_putreg27_in[147:140], zll_main_putreg27_in[139:0]};
  assign zll_main_putreg1_in = {zll_main_putreg_in[147:140], zll_main_putreg_in[139:70]};
  assign res = {zll_main_putreg1_in[77:70], zll_main_putreg1_in[61:54], zll_main_putreg1_in[53:46], zll_main_putreg1_in[45:38], zll_main_putreg1_in[37:32], zll_main_putreg1_in[31:15], zll_main_putreg1_in[14:0]};
endmodule

module ZLL_Main_r02 (input logic [7:0] arg0,
  input logic [5:0] arg1,
  input logic [16:0] arg2,
  input logic [14:0] arg3,
  output logic [7:0] res);
  logic [39:0] zll_main_r01_in;
  logic [22:0] zll_main_r0_in;
  assign zll_main_r01_in = {arg0, arg2, arg3};
  assign zll_main_r0_in = {zll_main_r01_in[39:32], zll_main_r01_in[14:0]};
  assign res = zll_main_r0_in[22:15];
endmodule

module ZLL_Main_r03 (input logic [7:0] arg0,
  input logic [7:0] arg1,
  input logic [5:0] arg2,
  input logic [16:0] arg3,
  input logic [14:0] arg4,
  output logic [7:0] res);
  logic [45:0] zll_main_r02_in;
  logic [7:0] zll_main_r02_out;
  assign zll_main_r02_in = {arg0, arg2, arg3, arg4};
  ZLL_Main_r02  inst (zll_main_r02_in[45:38], zll_main_r02_in[37:32], zll_main_r02_in[31:15], zll_main_r02_in[14:0], zll_main_r02_out);
  assign res = zll_main_r02_out;
endmodule

module ZLL_Main_r04 (input logic [7:0] arg0,
  input logic [7:0] arg1,
  input logic [7:0] arg2,
  input logic [5:0] arg3,
  input logic [16:0] arg4,
  input logic [14:0] arg5,
  output logic [7:0] res);
  logic [53:0] zll_main_r03_in;
  logic [7:0] zll_main_r03_out;
  assign zll_main_r03_in = {arg0, arg2, arg3, arg4, arg5};
  ZLL_Main_r03  inst (zll_main_r03_in[53:46], zll_main_r03_in[45:38], zll_main_r03_in[37:32], zll_main_r03_in[31:15], zll_main_r03_in[14:0], zll_main_r03_out);
  assign res = zll_main_r03_out;
endmodule

module ZLL_Pure_dispatch2 (input logic [16:0] arg0,
  input logic [69:0] arg1,
  output logic [142:0] res);
  logic [86:0] zll_main_loop1_in;
  logic [86:0] main_putins_in;
  logic [69:0] main_putins_out;
  logic [69:0] zll_main_loop87_in;
  logic [142:0] zll_main_loop87_out;
  logic [142:0] zll_main_loop86_in;
  logic [142:0] zll_main_loop86_out;
  assign zll_main_loop1_in = {arg0, arg1};
  assign main_putins_in = {zll_main_loop1_in[86:70], zll_main_loop1_in[69:0]};
  Main_putIns  inst (main_putins_in[86:70], main_putins_in[69:0], main_putins_out);
  assign zll_main_loop87_in = main_putins_out;
  ZLL_Main_loop87  instR1 (zll_main_loop87_in[69:0], zll_main_loop87_out);
  assign zll_main_loop86_in = zll_main_loop87_out;
  ZLL_Main_loop86  instR2 (zll_main_loop86_in[142:0], zll_main_loop86_out);
  assign res = zll_main_loop86_out;
endmodule

module Main_getIns (input logic [69:0] arg0,
  output logic [86:0] res);
  logic [139:0] zll_main_getins2_in;
  logic [139:0] zll_main_getins_in;
  logic [69:0] main_inputs_in;
  logic [69:0] zll_main_inputs6_in;
  logic [61:0] zll_main_inputs5_in;
  logic [53:0] zll_main_inputs4_in;
  logic [45:0] zll_main_inputs3_in;
  logic [37:0] zll_main_inputs2_in;
  logic [31:0] zll_main_inputs_in;
  assign zll_main_getins2_in = {arg0, arg0};
  assign zll_main_getins_in = zll_main_getins2_in[139:0];
  assign main_inputs_in = zll_main_getins_in[139:70];
  assign zll_main_inputs6_in = main_inputs_in[69:0];
  assign zll_main_inputs5_in = {zll_main_inputs6_in[61:54], zll_main_inputs6_in[53:46], zll_main_inputs6_in[45:38], zll_main_inputs6_in[37:32], zll_main_inputs6_in[31:15], zll_main_inputs6_in[14:0]};
  assign zll_main_inputs4_in = {zll_main_inputs5_in[53:46], zll_main_inputs5_in[45:38], zll_main_inputs5_in[37:32], zll_main_inputs5_in[31:15], zll_main_inputs5_in[14:0]};
  assign zll_main_inputs3_in = {zll_main_inputs4_in[45:38], zll_main_inputs4_in[37:32], zll_main_inputs4_in[31:15], zll_main_inputs4_in[14:0]};
  assign zll_main_inputs2_in = {zll_main_inputs3_in[37:32], zll_main_inputs3_in[31:15], zll_main_inputs3_in[14:0]};
  assign zll_main_inputs_in = {zll_main_inputs2_in[31:15], zll_main_inputs2_in[14:0]};
  assign res = {zll_main_inputs_in[31:15], zll_main_getins_in[69:0]};
endmodule

module Main_getOut (input logic [69:0] arg0,
  output logic [84:0] res);
  logic [139:0] zll_main_getout2_in;
  logic [139:0] zll_main_getout_in;
  logic [69:0] main_outputs_in;
  logic [69:0] zll_main_outputs6_in;
  logic [61:0] zll_main_outputs5_in;
  logic [53:0] zll_main_outputs4_in;
  logic [45:0] zll_main_outputs3_in;
  logic [37:0] zll_main_outputs2_in;
  logic [31:0] zll_main_outputs1_in;
  assign zll_main_getout2_in = {arg0, arg0};
  assign zll_main_getout_in = zll_main_getout2_in[139:0];
  assign main_outputs_in = zll_main_getout_in[139:70];
  assign zll_main_outputs6_in = main_outputs_in[69:0];
  assign zll_main_outputs5_in = {zll_main_outputs6_in[61:54], zll_main_outputs6_in[53:46], zll_main_outputs6_in[45:38], zll_main_outputs6_in[37:32], zll_main_outputs6_in[31:15], zll_main_outputs6_in[14:0]};
  assign zll_main_outputs4_in = {zll_main_outputs5_in[53:46], zll_main_outputs5_in[45:38], zll_main_outputs5_in[37:32], zll_main_outputs5_in[31:15], zll_main_outputs5_in[14:0]};
  assign zll_main_outputs3_in = {zll_main_outputs4_in[45:38], zll_main_outputs4_in[37:32], zll_main_outputs4_in[31:15], zll_main_outputs4_in[14:0]};
  assign zll_main_outputs2_in = {zll_main_outputs3_in[37:32], zll_main_outputs3_in[31:15], zll_main_outputs3_in[14:0]};
  assign zll_main_outputs1_in = {zll_main_outputs2_in[31:15], zll_main_outputs2_in[14:0]};
  assign res = {zll_main_outputs1_in[14:0], zll_main_getout_in[69:0]};
endmodule

module Main_getPC (input logic [69:0] arg0,
  output logic [75:0] res);
  logic [139:0] zll_main_getpc2_in;
  logic [139:0] zll_main_getpc_in;
  logic [69:0] main_pc_in;
  logic [69:0] zll_main_pc6_in;
  logic [61:0] zll_main_pc5_in;
  logic [53:0] zll_main_pc4_in;
  logic [45:0] zll_main_pc3_in;
  logic [37:0] zll_main_pc1_in;
  logic [20:0] zll_main_pc_in;
  assign zll_main_getpc2_in = {arg0, arg0};
  assign zll_main_getpc_in = zll_main_getpc2_in[139:0];
  assign main_pc_in = zll_main_getpc_in[139:70];
  assign zll_main_pc6_in = main_pc_in[69:0];
  assign zll_main_pc5_in = {zll_main_pc6_in[61:54], zll_main_pc6_in[53:46], zll_main_pc6_in[45:38], zll_main_pc6_in[37:32], zll_main_pc6_in[31:15], zll_main_pc6_in[14:0]};
  assign zll_main_pc4_in = {zll_main_pc5_in[53:46], zll_main_pc5_in[45:38], zll_main_pc5_in[37:32], zll_main_pc5_in[31:15], zll_main_pc5_in[14:0]};
  assign zll_main_pc3_in = {zll_main_pc4_in[45:38], zll_main_pc4_in[37:32], zll_main_pc4_in[31:15], zll_main_pc4_in[14:0]};
  assign zll_main_pc1_in = {zll_main_pc3_in[37:32], zll_main_pc3_in[31:15], zll_main_pc3_in[14:0]};
  assign zll_main_pc_in = {zll_main_pc1_in[37:32], zll_main_pc1_in[14:0]};
  assign res = {zll_main_pc_in[20:15], zll_main_getpc_in[69:0]};
endmodule

module Main_getReg (input logic [1:0] arg0,
  input logic [69:0] arg1,
  output logic [77:0] res);
  logic [71:0] zll_main_getreg20_in;
  logic [69:0] zll_main_getreg8_in;
  logic [139:0] zll_main_getreg16_in;
  logic [139:0] zll_main_getreg3_in;
  logic [69:0] main_r3_in;
  logic [69:0] zll_main_r36_in;
  logic [61:0] zll_main_r35_in;
  logic [53:0] zll_main_r34_in;
  logic [45:0] zll_main_r02_in;
  logic [7:0] zll_main_r02_out;
  logic [71:0] zll_main_getreg19_in;
  logic [69:0] zll_main_getreg7_in;
  logic [139:0] zll_main_getreg14_in;
  logic [139:0] zll_main_getreg2_in;
  logic [69:0] main_r2_in;
  logic [69:0] zll_main_r26_in;
  logic [61:0] zll_main_r25_in;
  logic [53:0] zll_main_r03_in;
  logic [7:0] zll_main_r03_out;
  logic [71:0] zll_main_getreg18_in;
  logic [69:0] zll_main_getreg6_in;
  logic [139:0] zll_main_getreg12_in;
  logic [139:0] zll_main_getreg1_in;
  logic [69:0] main_r1_in;
  logic [69:0] zll_main_r16_in;
  logic [61:0] zll_main_r04_in;
  logic [7:0] zll_main_r04_out;
  logic [71:0] zll_main_getreg17_in;
  logic [69:0] zll_main_getreg5_in;
  logic [77:0] zll_main_getreg5_out;
  assign zll_main_getreg20_in = {arg1, arg0};
  assign zll_main_getreg8_in = zll_main_getreg20_in[71:2];
  assign zll_main_getreg16_in = {zll_main_getreg8_in[69:0], zll_main_getreg8_in[69:0]};
  assign zll_main_getreg3_in = zll_main_getreg16_in[139:0];
  assign main_r3_in = zll_main_getreg3_in[139:70];
  assign zll_main_r36_in = main_r3_in[69:0];
  assign zll_main_r35_in = {zll_main_r36_in[61:54], zll_main_r36_in[53:46], zll_main_r36_in[45:38], zll_main_r36_in[37:32], zll_main_r36_in[31:15], zll_main_r36_in[14:0]};
  assign zll_main_r34_in = {zll_main_r35_in[53:46], zll_main_r35_in[45:38], zll_main_r35_in[37:32], zll_main_r35_in[31:15], zll_main_r35_in[14:0]};
  assign zll_main_r02_in = {zll_main_r34_in[45:38], zll_main_r34_in[37:32], zll_main_r34_in[31:15], zll_main_r34_in[14:0]};
  ZLL_Main_r02  inst (zll_main_r02_in[45:38], zll_main_r02_in[37:32], zll_main_r02_in[31:15], zll_main_r02_in[14:0], zll_main_r02_out);
  assign zll_main_getreg19_in = {arg1, arg0};
  assign zll_main_getreg7_in = zll_main_getreg19_in[71:2];
  assign zll_main_getreg14_in = {zll_main_getreg7_in[69:0], zll_main_getreg7_in[69:0]};
  assign zll_main_getreg2_in = zll_main_getreg14_in[139:0];
  assign main_r2_in = zll_main_getreg2_in[139:70];
  assign zll_main_r26_in = main_r2_in[69:0];
  assign zll_main_r25_in = {zll_main_r26_in[61:54], zll_main_r26_in[53:46], zll_main_r26_in[45:38], zll_main_r26_in[37:32], zll_main_r26_in[31:15], zll_main_r26_in[14:0]};
  assign zll_main_r03_in = {zll_main_r25_in[53:46], zll_main_r25_in[45:38], zll_main_r25_in[37:32], zll_main_r25_in[31:15], zll_main_r25_in[14:0]};
  ZLL_Main_r03  instR1 (zll_main_r03_in[53:46], zll_main_r03_in[45:38], zll_main_r03_in[37:32], zll_main_r03_in[31:15], zll_main_r03_in[14:0], zll_main_r03_out);
  assign zll_main_getreg18_in = {arg1, arg0};
  assign zll_main_getreg6_in = zll_main_getreg18_in[71:2];
  assign zll_main_getreg12_in = {zll_main_getreg6_in[69:0], zll_main_getreg6_in[69:0]};
  assign zll_main_getreg1_in = zll_main_getreg12_in[139:0];
  assign main_r1_in = zll_main_getreg1_in[139:70];
  assign zll_main_r16_in = main_r1_in[69:0];
  assign zll_main_r04_in = {zll_main_r16_in[61:54], zll_main_r16_in[53:46], zll_main_r16_in[45:38], zll_main_r16_in[37:32], zll_main_r16_in[31:15], zll_main_r16_in[14:0]};
  ZLL_Main_r04  instR2 (zll_main_r04_in[61:54], zll_main_r04_in[53:46], zll_main_r04_in[45:38], zll_main_r04_in[37:32], zll_main_r04_in[31:15], zll_main_r04_in[14:0], zll_main_r04_out);
  assign zll_main_getreg17_in = {arg1, arg0};
  assign zll_main_getreg5_in = zll_main_getreg17_in[71:2];
  ZLL_Main_getReg5  instR3 (zll_main_getreg5_in[69:0], zll_main_getreg5_out);
  assign res = (zll_main_getreg17_in[1:0] == 2'h0) ? zll_main_getreg5_out : ((zll_main_getreg18_in[1:0] == 2'h1) ? {zll_main_r04_out, zll_main_getreg1_in[69:0]} : ((zll_main_getreg19_in[1:0] == 2'h2) ? {zll_main_r03_out, zll_main_getreg2_in[69:0]} : {zll_main_r02_out, zll_main_getreg3_in[69:0]}));
endmodule

module Main_incrPC (input logic [69:0] arg0,
  output logic [69:0] res);
  logic [69:0] main_getpc_in;
  logic [75:0] main_getpc_out;
  logic [75:0] zll_main_incrpc2_in;
  logic [75:0] zll_main_incrpc_in;
  logic [11:0] binop_in;
  logic [75:0] main_putpc_in;
  logic [69:0] main_putpc_out;
  assign main_getpc_in = arg0;
  Main_getPC  inst (main_getpc_in[69:0], main_getpc_out);
  assign zll_main_incrpc2_in = main_getpc_out;
  assign zll_main_incrpc_in = zll_main_incrpc2_in[75:0];
  assign binop_in = {zll_main_incrpc_in[75:70], 6'h01};
  assign main_putpc_in = {binop_in[11:6] + binop_in[5:0], zll_main_incrpc_in[69:0]};
  Main_putPC  instR1 (main_putpc_in[75:70], main_putpc_in[69:0], main_putpc_out);
  assign res = main_putpc_out;
endmodule

module Main_putAddrOut (input logic [5:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [69:0] main_getout_in;
  logic [84:0] main_getout_out;
  logic [90:0] zll_main_putaddrout6_in;
  logic [90:0] zll_main_putaddrout_in;
  logic [20:0] zll_main_putaddrout1_in;
  logic [84:0] main_putout_in;
  logic [69:0] main_putout_out;
  assign main_getout_in = arg1;
  Main_getOut  inst (main_getout_in[69:0], main_getout_out);
  assign zll_main_putaddrout6_in = {arg0, main_getout_out};
  assign zll_main_putaddrout_in = {zll_main_putaddrout6_in[90:85], zll_main_putaddrout6_in[84:0]};
  assign zll_main_putaddrout1_in = {zll_main_putaddrout_in[90:85], zll_main_putaddrout_in[84:70]};
  assign main_putout_in = {{zll_main_putaddrout1_in[14], zll_main_putaddrout1_in[20:15], zll_main_putaddrout1_in[7:0]}, zll_main_putaddrout_in[69:0]};
  Main_putOut  instR1 (main_putout_in[84:70], main_putout_in[69:0], main_putout_out);
  assign res = main_putout_out;
endmodule

module Main_putIns (input logic [16:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [156:0] zll_main_putins10_in;
  logic [156:0] zll_main_putins_in;
  logic [86:0] zll_main_putins6_in;
  logic [86:0] zll_main_putins5_in;
  logic [86:0] zll_main_putins4_in;
  logic [86:0] zll_main_putins2_in;
  logic [86:0] zll_main_putins1_in;
  assign zll_main_putins10_in = {arg0, arg1, arg1};
  assign zll_main_putins_in = {zll_main_putins10_in[156:140], zll_main_putins10_in[139:0]};
  assign zll_main_putins6_in = {zll_main_putins_in[156:140], zll_main_putins_in[139:70]};
  assign zll_main_putins5_in = {zll_main_putins6_in[69:62], zll_main_putins6_in[86:70], zll_main_putins6_in[61:54], zll_main_putins6_in[53:46], zll_main_putins6_in[45:38], zll_main_putins6_in[37:32], zll_main_putins6_in[31:15], zll_main_putins6_in[14:0]};
  assign zll_main_putins4_in = {zll_main_putins5_in[61:54], zll_main_putins5_in[86:79], zll_main_putins5_in[78:62], zll_main_putins5_in[53:46], zll_main_putins5_in[45:38], zll_main_putins5_in[37:32], zll_main_putins5_in[31:15], zll_main_putins5_in[14:0]};
  assign zll_main_putins2_in = {zll_main_putins4_in[53:46], zll_main_putins4_in[86:79], zll_main_putins4_in[78:71], zll_main_putins4_in[70:54], zll_main_putins4_in[45:38], zll_main_putins4_in[37:32], zll_main_putins4_in[31:15], zll_main_putins4_in[14:0]};
  assign zll_main_putins1_in = {zll_main_putins2_in[86:79], zll_main_putins2_in[78:71], zll_main_putins2_in[70:63], zll_main_putins2_in[37:32], zll_main_putins2_in[62:46], zll_main_putins2_in[45:38], zll_main_putins2_in[31:15], zll_main_putins2_in[14:0]};
  assign res = {zll_main_putins1_in[70:63], zll_main_putins1_in[78:71], zll_main_putins1_in[86:79], zll_main_putins1_in[39:32], zll_main_putins1_in[62:57], zll_main_putins1_in[56:40], zll_main_putins1_in[14:0]};
endmodule

module Main_putOut (input logic [14:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [154:0] zll_main_putout11_in;
  logic [154:0] zll_main_putout_in;
  logic [84:0] zll_main_putout7_in;
  logic [84:0] zll_main_putout6_in;
  logic [84:0] zll_main_putout4_in;
  logic [84:0] zll_main_putout3_in;
  logic [84:0] zll_main_putout2_in;
  logic [84:0] zll_main_putout1_in;
  assign zll_main_putout11_in = {arg0, arg1, arg1};
  assign zll_main_putout_in = {zll_main_putout11_in[154:140], zll_main_putout11_in[139:0]};
  assign zll_main_putout7_in = {zll_main_putout_in[154:140], zll_main_putout_in[139:70]};
  assign zll_main_putout6_in = {zll_main_putout7_in[69:62], zll_main_putout7_in[84:70], zll_main_putout7_in[61:54], zll_main_putout7_in[53:46], zll_main_putout7_in[45:38], zll_main_putout7_in[37:32], zll_main_putout7_in[31:15], zll_main_putout7_in[14:0]};
  assign zll_main_putout4_in = {zll_main_putout6_in[61:54], zll_main_putout6_in[84:77], zll_main_putout6_in[76:62], zll_main_putout6_in[53:46], zll_main_putout6_in[45:38], zll_main_putout6_in[37:32], zll_main_putout6_in[31:15], zll_main_putout6_in[14:0]};
  assign zll_main_putout3_in = {zll_main_putout4_in[45:38], zll_main_putout4_in[84:77], zll_main_putout4_in[76:69], zll_main_putout4_in[68:54], zll_main_putout4_in[53:46], zll_main_putout4_in[37:32], zll_main_putout4_in[31:15], zll_main_putout4_in[14:0]};
  assign zll_main_putout2_in = {zll_main_putout3_in[37:32], zll_main_putout3_in[84:77], zll_main_putout3_in[76:69], zll_main_putout3_in[68:61], zll_main_putout3_in[60:46], zll_main_putout3_in[45:38], zll_main_putout3_in[31:15], zll_main_putout3_in[14:0]};
  assign zll_main_putout1_in = {zll_main_putout2_in[84:79], zll_main_putout2_in[78:71], zll_main_putout2_in[70:63], zll_main_putout2_in[62:55], zll_main_putout2_in[54:40], zll_main_putout2_in[31:15], zll_main_putout2_in[39:32], zll_main_putout2_in[14:0]};
  assign res = {zll_main_putout1_in[62:55], zll_main_putout1_in[70:63], zll_main_putout1_in[22:15], zll_main_putout1_in[78:71], zll_main_putout1_in[84:79], zll_main_putout1_in[39:23], zll_main_putout1_in[54:40]};
endmodule

module Main_putPC (input logic [5:0] arg0,
  input logic [69:0] arg1,
  output logic [69:0] res);
  logic [145:0] zll_main_putpc15_in;
  logic [145:0] zll_main_putpc_in;
  logic [75:0] zll_main_putpc4_in;
  logic [75:0] zll_main_putpc3_in;
  logic [75:0] zll_main_putpc2_in;
  logic [75:0] zll_main_putpc1_in;
  assign zll_main_putpc15_in = {arg0, arg1, arg1};
  assign zll_main_putpc_in = {zll_main_putpc15_in[145:140], zll_main_putpc15_in[139:0]};
  assign zll_main_putpc4_in = {zll_main_putpc_in[145:140], zll_main_putpc_in[139:70]};
  assign zll_main_putpc3_in = {zll_main_putpc4_in[61:54], zll_main_putpc4_in[75:70], zll_main_putpc4_in[69:62], zll_main_putpc4_in[53:46], zll_main_putpc4_in[45:38], zll_main_putpc4_in[37:32], zll_main_putpc4_in[31:15], zll_main_putpc4_in[14:0]};
  assign zll_main_putpc2_in = {zll_main_putpc3_in[53:46], zll_main_putpc3_in[75:68], zll_main_putpc3_in[67:62], zll_main_putpc3_in[61:54], zll_main_putpc3_in[45:38], zll_main_putpc3_in[37:32], zll_main_putpc3_in[31:15], zll_main_putpc3_in[14:0]};
  assign zll_main_putpc1_in = {zll_main_putpc2_in[75:68], zll_main_putpc2_in[45:38], zll_main_putpc2_in[67:60], zll_main_putpc2_in[59:54], zll_main_putpc2_in[53:46], zll_main_putpc2_in[37:32], zll_main_putpc2_in[31:15], zll_main_putpc2_in[14:0]};
  assign res = {zll_main_putpc1_in[45:38], zll_main_putpc1_in[59:52], zll_main_putpc1_in[75:68], zll_main_putpc1_in[67:60], zll_main_putpc1_in[51:46], zll_main_putpc1_in[31:15], zll_main_putpc1_in[14:0]};
endmodule

module Main_putWeOut (input logic [69:0] arg0,
  output logic [69:0] res);
  logic [69:0] main_getout_in;
  logic [84:0] main_getout_out;
  logic [84:0] zll_main_putweout5_in;
  logic [84:0] zll_main_putweout_in;
  logic [14:0] zll_main_putweout1_in;
  logic [84:0] main_putout_in;
  logic [69:0] main_putout_out;
  assign main_getout_in = arg0;
  Main_getOut  inst (main_getout_in[69:0], main_getout_out);
  assign zll_main_putweout5_in = main_getout_out;
  assign zll_main_putweout_in = zll_main_putweout5_in[84:0];
  assign zll_main_putweout1_in = zll_main_putweout_in[84:70];
  assign main_putout_in = {{1'h0, zll_main_putweout1_in[13:8], zll_main_putweout1_in[7:0]}, zll_main_putweout_in[69:0]};
  Main_putOut  instR1 (main_putout_in[84:70], main_putout_in[69:0], main_putout_out);
  assign res = main_putout_out;
endmodule