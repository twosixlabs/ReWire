module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [9:0] __in0,
  output logic [15:0] __out0);
  logic [39:0] rewire_monad_iterst1_in;
  logic [69:0] zll_rewire_monad_iterst42_in;
  logic [69:0] zll_rewire_monad_iterst9_in;
  logic [39:0] main_loop_in;
  logic [29:0] id_in;
  logic [24:0] main_inputtomystate_in;
  logic [24:0] zll_main_inputtomystate13_in;
  logic [13:0] zll_main_inputtomystate12_in;
  logic [24:0] zll_main_inputtomystate11_in;
  logic [24:0] zll_main_inputtomystate10_in;
  logic [12:0] zll_main_inputtomystate8_in;
  logic [24:0] zll_main_inputtomystate6_in;
  logic [22:0] zll_main_inputtomystate5_in;
  logic [22:0] zll_main_inputtomystate4_in;
  logic [24:0] zll_main_inputtomystate2_in;
  logic [18:0] zll_main_inputtomystate1_in;
  logic [13:0] zll_main_inputtomystate_in;
  logic [44:0] main_incrpipeline_in;
  logic [44:0] zll_main_incrpipeline_in;
  logic [29:0] id_inR1;
  logic [29:0] resize_in;
  logic [255:0] binop_in;
  logic [127:0] resize_inR1;
  logic [44:0] zll_main_loop_in;
  logic [14:0] main_mystatetooutput_in;
  logic [14:0] zll_main_mystatetooutput5_in;
  logic [8:0] zll_main_mystatetooutput4_in;
  logic [14:0] zll_main_mystatetooutput3_in;
  logic [12:0] zll_main_mystatetooutput2_in;
  logic [14:0] zll_main_mystatetooutput1_in;
  logic [8:0] zll_main_mystatetooutput_in;
  logic [75:0] zll_rewire_monad_iterst39_in;
  logic [75:0] zll_rewire_monad_iterst30_in;
  logic [77:0] zll_rewire_monad_iterst36_in;
  logic [77:0] zll_rewire_monad_iterst35_in;
  logic [75:0] zll_rewire_monad_iterst6_in;
  logic [75:0] zll_rewire_monad_iterst20_in;
  logic [75:0] zll_rewire_monad_iterst19_in;
  logic [75:0] zll_rewire_monad_iterst7_in;
  logic [29:0] zll_rewire_monad_iterst16_in;
  logic [93:0] zll_rewire_monad_iterst24_in;
  logic [93:0] zll_rewire_monad_iterst22_in;
  logic [45:0] zll_rewire_monad_iterst_in;
  logic [0:0] __continue;
  logic [30:0] __padding;
  logic [29:0] __st0;
  logic [29:0] __st0_next;
  assign rewire_monad_iterst1_in = {__in0, __st0};
  assign zll_rewire_monad_iterst42_in = {rewire_monad_iterst1_in[39:30], rewire_monad_iterst1_in[29:0], rewire_monad_iterst1_in[29:0]};
  assign zll_rewire_monad_iterst9_in = {zll_rewire_monad_iterst42_in[69:60], zll_rewire_monad_iterst42_in[59:0]};
  assign main_loop_in = {zll_rewire_monad_iterst9_in[69:60], zll_rewire_monad_iterst9_in[59:30]};
  assign id_in = main_loop_in[29:0];
  assign main_inputtomystate_in = {main_loop_in[39:30], id_in[29:15]};
  assign zll_main_inputtomystate13_in = {main_inputtomystate_in[24:15], main_inputtomystate_in[14:0]};
  assign zll_main_inputtomystate12_in = {zll_main_inputtomystate13_in[13:9], zll_main_inputtomystate13_in[8:0]};
  assign zll_main_inputtomystate11_in = {main_inputtomystate_in[24:15], main_inputtomystate_in[14:0]};
  assign zll_main_inputtomystate10_in = {main_inputtomystate_in[24:15], main_inputtomystate_in[14:0]};
  assign zll_main_inputtomystate8_in = {zll_main_inputtomystate10_in[12:9], zll_main_inputtomystate10_in[8:0]};
  assign zll_main_inputtomystate6_in = {main_inputtomystate_in[24:15], main_inputtomystate_in[14:0]};
  assign zll_main_inputtomystate5_in = {zll_main_inputtomystate6_in[22:15], zll_main_inputtomystate6_in[14], zll_main_inputtomystate6_in[13:9], zll_main_inputtomystate6_in[8:0]};
  assign zll_main_inputtomystate4_in = {zll_main_inputtomystate5_in[22:15], zll_main_inputtomystate5_in[13:9], zll_main_inputtomystate5_in[14], zll_main_inputtomystate5_in[8:0]};
  assign zll_main_inputtomystate2_in = {main_inputtomystate_in[24:15], main_inputtomystate_in[14:0]};
  assign zll_main_inputtomystate1_in = {zll_main_inputtomystate2_in[18:15], zll_main_inputtomystate2_in[14], zll_main_inputtomystate2_in[13:9], zll_main_inputtomystate2_in[8:0]};
  assign zll_main_inputtomystate_in = {zll_main_inputtomystate1_in[18:15], zll_main_inputtomystate1_in[14], zll_main_inputtomystate1_in[8:0]};
  assign main_incrpipeline_in = {(zll_main_inputtomystate2_in[24:23] == 2'h0) ? {zll_main_inputtomystate_in[9], 1'h1, zll_main_inputtomystate_in[13:10], 5'h00, zll_main_inputtomystate_in[13:10]} : ((zll_main_inputtomystate6_in[24:23] == 2'h1) ? {zll_main_inputtomystate4_in[9], zll_main_inputtomystate4_in[14:10], 1'h1, zll_main_inputtomystate4_in[22:15]} : (((zll_main_inputtomystate10_in[24:23] == 2'h2) && ((zll_main_inputtomystate10_in[15] == 1'h1) && (zll_main_inputtomystate10_in[13] == 1'h1))) ? {11'h400, zll_main_inputtomystate8_in[12:9]} : (((zll_main_inputtomystate11_in[24:23] == 2'h2) && ((zll_main_inputtomystate11_in[15] == 1'h1) && (zll_main_inputtomystate11_in[13] == 1'h0))) ? {6'h20, zll_main_inputtomystate11_in[8:0]} : {6'h00, zll_main_inputtomystate12_in[8:0]}))), main_loop_in[29:0]};
  assign zll_main_incrpipeline_in = main_incrpipeline_in[44:0];
  assign id_inR1 = zll_main_incrpipeline_in[29:0];
  assign resize_in = zll_main_incrpipeline_in[29:0];
  assign binop_in = {128'(resize_in[29:0]), {8'h80{1'h0}}};
  assign resize_inR1 = binop_in[255:128] >> binop_in[127:0];
  assign zll_main_loop_in = {zll_main_incrpipeline_in[44:30], id_inR1[29:15], resize_inR1[14:0]};
  assign main_mystatetooutput_in = zll_main_loop_in[14:0];
  assign zll_main_mystatetooutput5_in = main_mystatetooutput_in[14:0];
  assign zll_main_mystatetooutput4_in = zll_main_mystatetooutput5_in[8:0];
  assign zll_main_mystatetooutput3_in = main_mystatetooutput_in[14:0];
  assign zll_main_mystatetooutput2_in = {zll_main_mystatetooutput3_in[13:9], zll_main_mystatetooutput3_in[7:0]};
  assign zll_main_mystatetooutput1_in = main_mystatetooutput_in[14:0];
  assign zll_main_mystatetooutput_in = {zll_main_mystatetooutput1_in[13:9], zll_main_mystatetooutput1_in[3:0]};
  assign zll_rewire_monad_iterst39_in = {{((zll_main_mystatetooutput1_in[14] == 1'h1) && (zll_main_mystatetooutput1_in[8] == 1'h0)) ? {2'h3, zll_main_mystatetooutput_in[8:4], 5'h00, zll_main_mystatetooutput_in[3:0]} : (((zll_main_mystatetooutput3_in[14] == 1'h1) && (zll_main_mystatetooutput3_in[8] == 1'h1)) ? {2'h1, zll_main_mystatetooutput2_in[12:8], 1'h1, zll_main_mystatetooutput2_in[7:0]} : {7'h00, zll_main_mystatetooutput4_in[8:0]}), zll_main_loop_in[44:15]}, zll_rewire_monad_iterst9_in[29:0]};
  assign zll_rewire_monad_iterst30_in = zll_rewire_monad_iterst39_in[75:0];
  assign zll_rewire_monad_iterst36_in = {2'h0, zll_rewire_monad_iterst30_in[75:30], zll_rewire_monad_iterst30_in[29:0]};
  assign zll_rewire_monad_iterst35_in = zll_rewire_monad_iterst36_in[77:0];
  assign zll_rewire_monad_iterst6_in = {zll_rewire_monad_iterst35_in[75:30], zll_rewire_monad_iterst35_in[29:0]};
  assign zll_rewire_monad_iterst20_in = {zll_rewire_monad_iterst6_in[29:0], zll_rewire_monad_iterst6_in[75:30]};
  assign zll_rewire_monad_iterst19_in = {zll_rewire_monad_iterst20_in[45:30], zll_rewire_monad_iterst20_in[75:46], zll_rewire_monad_iterst20_in[29:0]};
  assign zll_rewire_monad_iterst7_in = {zll_rewire_monad_iterst19_in[75:60], zll_rewire_monad_iterst19_in[29:0], zll_rewire_monad_iterst19_in[59:30]};
  assign zll_rewire_monad_iterst16_in = zll_rewire_monad_iterst7_in[59:30];
  assign zll_rewire_monad_iterst24_in = {zll_rewire_monad_iterst7_in[75:60], {{2'h1, {6'h2e{1'h0}}}, zll_rewire_monad_iterst16_in[29:0]}};
  assign zll_rewire_monad_iterst22_in = {zll_rewire_monad_iterst24_in[93:78], zll_rewire_monad_iterst24_in[77:0]};
  assign zll_rewire_monad_iterst_in = {zll_rewire_monad_iterst22_in[93:78], zll_rewire_monad_iterst22_in[29:0]};
  assign {__continue, __padding, __out0, __st0_next} = {{1'h1, {5'h1f{1'h0}}}, zll_rewire_monad_iterst_in[45:30], zll_rewire_monad_iterst_in[29:0]};
  initial __st0 <= 30'h00000000;
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      __st0 <= 30'h00000000;
    end else begin
      __st0 <= __st0_next;
    end
  end
endmodule