module top_level (input logic [7:0] __in0,
  output logic [7:0] __out0,
  output logic [7:0] __out1,
  output logic [7:0] __out2,
  output logic [7:0] __out3);
  logic [7:0] zll_main_dev226_in;
  logic [7:0] zll_main_x2_in;
  logic [15:0] binop_in;
  logic [15:0] zll_main_dev136_in;
  logic [15:0] zll_main_dev22_in;
  logic [15:0] zll_main_dev233_in;
  logic [15:0] zll_main_dev239_in;
  logic [15:0] zll_main_dev19_in;
  logic [18:0] zll_main_dev128_in;
  logic [18:0] zll_main_dev261_in;
  logic [21:0] zll_main_dev84_in;
  logic [24:0] zll_main_dev18_in;
  logic [0:0] zll_main_dev18_out;
  logic [24:0] zll_main_dev18_inR1;
  logic [0:0] zll_main_dev18_outR1;
  logic [24:0] zll_main_dev18_inR2;
  logic [0:0] zll_main_dev18_outR2;
  logic [24:0] zll_main_dev18_inR3;
  logic [0:0] zll_main_dev18_outR3;
  logic [24:0] zll_main_dev18_inR4;
  logic [0:0] zll_main_dev18_outR4;
  logic [24:0] zll_main_dev18_inR5;
  logic [0:0] zll_main_dev18_outR5;
  logic [24:0] zll_main_dev18_inR6;
  logic [0:0] zll_main_dev18_outR6;
  logic [24:0] zll_main_dev18_inR7;
  logic [0:0] zll_main_dev18_outR7;
  logic [15:0] zll_main_dev250_in;
  logic [15:0] zll_main_dev253_in;
  logic [15:0] zll_main_dev17_in;
  logic [15:0] zll_main_dev197_in;
  logic [18:0] zll_main_dev3_in;
  logic [21:0] zll_main_dev69_in;
  logic [5:0] zll_main_dev262_in;
  logic [2:0] zll_main_dev262_out;
  logic [24:0] zll_main_dev252_in;
  logic [14:0] zll_main_dev87_in;
  logic [6:0] zll_main_dev176_in;
  logic [2:0] zll_main_dev176_out;
  logic [3:0] id_in;
  logic [24:0] zll_main_dev5_in;
  logic [27:0] zll_main_dev221_in;
  logic [0:0] zll_main_dev221_out;
  logic [27:0] zll_main_dev221_inR1;
  logic [0:0] zll_main_dev221_outR1;
  logic [27:0] zll_main_dev221_inR2;
  logic [0:0] zll_main_dev221_outR2;
  logic [27:0] zll_main_dev221_inR3;
  logic [0:0] zll_main_dev221_outR3;
  logic [27:0] zll_main_dev221_inR4;
  logic [0:0] zll_main_dev221_outR4;
  logic [27:0] zll_main_dev221_inR5;
  logic [0:0] zll_main_dev221_outR5;
  logic [27:0] zll_main_dev221_inR6;
  logic [0:0] zll_main_dev221_outR6;
  logic [27:0] zll_main_dev221_inR7;
  logic [0:0] zll_main_dev221_outR7;
  logic [15:0] zll_main_dev142_in;
  logic [15:0] zll_main_dev245_in;
  logic [15:0] zll_main_dev99_in;
  logic [15:0] zll_main_dev120_in;
  logic [18:0] zll_main_dev74_in;
  logic [18:0] zll_main_dev215_in;
  logic [21:0] zll_main_dev218_in;
  logic [5:0] zll_main_dev262_inR1;
  logic [2:0] zll_main_dev262_outR1;
  logic [24:0] zll_main_dev125_in;
  logic [14:0] zll_main_dev205_in;
  logic [6:0] zll_main_dev103_in;
  logic [6:0] zll_main_dev285_in;
  logic [5:0] zll_main_dev270_in;
  logic [2:0] zll_main_dev270_out;
  logic [3:0] id_inR1;
  logic [21:0] zll_main_dev202_in;
  logic [24:0] zll_main_dev101_in;
  logic [0:0] zll_main_dev101_out;
  logic [24:0] zll_main_dev101_inR1;
  logic [0:0] zll_main_dev101_outR1;
  logic [24:0] zll_main_dev101_inR2;
  logic [0:0] zll_main_dev101_outR2;
  logic [24:0] zll_main_dev101_inR3;
  logic [0:0] zll_main_dev101_outR3;
  logic [24:0] zll_main_dev101_inR4;
  logic [0:0] zll_main_dev101_outR4;
  logic [24:0] zll_main_dev101_inR5;
  logic [0:0] zll_main_dev101_outR5;
  logic [24:0] zll_main_dev101_inR6;
  logic [0:0] zll_main_dev101_outR6;
  logic [24:0] zll_main_dev101_inR7;
  logic [0:0] zll_main_dev101_outR7;
  logic [15:0] zll_main_dev234_in;
  logic [15:0] zll_main_dev38_in;
  logic [15:0] zll_main_dev169_in;
  logic [18:0] zll_main_dev37_in;
  logic [21:0] zll_main_dev42_in;
  logic [5:0] zll_main_dev262_inR2;
  logic [2:0] zll_main_dev262_outR2;
  logic [24:0] zll_main_dev171_in;
  logic [14:0] zll_main_dev89_in;
  logic [6:0] zll_main_dev176_inR1;
  logic [2:0] zll_main_dev176_outR1;
  logic [3:0] id_inR2;
  logic [24:0] zll_main_dev27_in;
  logic [27:0] zll_main_dev272_in;
  logic [0:0] zll_main_dev272_out;
  logic [27:0] zll_main_dev272_inR1;
  logic [0:0] zll_main_dev272_outR1;
  logic [27:0] zll_main_dev272_inR2;
  logic [0:0] zll_main_dev272_outR2;
  logic [27:0] zll_main_dev272_inR3;
  logic [0:0] zll_main_dev272_outR3;
  logic [27:0] zll_main_dev272_inR4;
  logic [0:0] zll_main_dev272_outR4;
  logic [27:0] zll_main_dev272_inR5;
  logic [0:0] zll_main_dev272_outR5;
  logic [27:0] zll_main_dev272_inR6;
  logic [0:0] zll_main_dev272_outR6;
  logic [27:0] zll_main_dev272_inR7;
  logic [0:0] zll_main_dev272_outR7;
  logic [0:0] __continue;
  assign zll_main_dev226_in = __in0;
  assign zll_main_x2_in = zll_main_dev226_in[7:0];
  assign binop_in = {zll_main_x2_in[7:0], 8'h2};
  assign zll_main_dev136_in = {zll_main_dev226_in[7:0], binop_in[15:8] * binop_in[7:0]};
  assign zll_main_dev22_in = {zll_main_dev136_in[15:8], zll_main_dev136_in[7:0]};
  assign zll_main_dev233_in = {zll_main_dev22_in[15:8], zll_main_dev22_in[7:0]};
  assign zll_main_dev239_in = zll_main_dev233_in[15:0];
  assign zll_main_dev19_in = {zll_main_dev239_in[7:0], zll_main_dev239_in[15:8]};
  assign zll_main_dev128_in = {zll_main_dev19_in[15:8], zll_main_dev19_in[7:0], 3'h1};
  assign zll_main_dev261_in = {zll_main_dev128_in[18:11], zll_main_dev128_in[2:0], zll_main_dev128_in[10:3]};
  assign zll_main_dev84_in = {zll_main_dev261_in[18:11], zll_main_dev261_in[10:8], zll_main_dev261_in[7:0], 3'h2};
  assign zll_main_dev18_in = {zll_main_dev84_in[2:0], zll_main_dev84_in[21:14], zll_main_dev84_in[13:11], zll_main_dev84_in[10:3], 3'h0};
  ZLL_Main_dev18  inst (zll_main_dev18_in[24:22], zll_main_dev18_in[21:14], zll_main_dev18_in[13:11], zll_main_dev18_in[10:3], zll_main_dev18_in[2:0], zll_main_dev18_out);
  assign zll_main_dev18_inR1 = {zll_main_dev84_in[2:0], zll_main_dev84_in[21:14], zll_main_dev84_in[13:11], zll_main_dev84_in[10:3], 3'h1};
  ZLL_Main_dev18  instR1 (zll_main_dev18_inR1[24:22], zll_main_dev18_inR1[21:14], zll_main_dev18_inR1[13:11], zll_main_dev18_inR1[10:3], zll_main_dev18_inR1[2:0], zll_main_dev18_outR1);
  assign zll_main_dev18_inR2 = {zll_main_dev84_in[2:0], zll_main_dev84_in[21:14], zll_main_dev84_in[13:11], zll_main_dev84_in[10:3], 3'h2};
  ZLL_Main_dev18  instR2 (zll_main_dev18_inR2[24:22], zll_main_dev18_inR2[21:14], zll_main_dev18_inR2[13:11], zll_main_dev18_inR2[10:3], zll_main_dev18_inR2[2:0], zll_main_dev18_outR2);
  assign zll_main_dev18_inR3 = {zll_main_dev84_in[2:0], zll_main_dev84_in[21:14], zll_main_dev84_in[13:11], zll_main_dev84_in[10:3], 3'h3};
  ZLL_Main_dev18  instR3 (zll_main_dev18_inR3[24:22], zll_main_dev18_inR3[21:14], zll_main_dev18_inR3[13:11], zll_main_dev18_inR3[10:3], zll_main_dev18_inR3[2:0], zll_main_dev18_outR3);
  assign zll_main_dev18_inR4 = {zll_main_dev84_in[2:0], zll_main_dev84_in[21:14], zll_main_dev84_in[13:11], zll_main_dev84_in[10:3], 3'h4};
  ZLL_Main_dev18  instR4 (zll_main_dev18_inR4[24:22], zll_main_dev18_inR4[21:14], zll_main_dev18_inR4[13:11], zll_main_dev18_inR4[10:3], zll_main_dev18_inR4[2:0], zll_main_dev18_outR4);
  assign zll_main_dev18_inR5 = {zll_main_dev84_in[2:0], zll_main_dev84_in[21:14], zll_main_dev84_in[13:11], zll_main_dev84_in[10:3], 3'h5};
  ZLL_Main_dev18  instR5 (zll_main_dev18_inR5[24:22], zll_main_dev18_inR5[21:14], zll_main_dev18_inR5[13:11], zll_main_dev18_inR5[10:3], zll_main_dev18_inR5[2:0], zll_main_dev18_outR5);
  assign zll_main_dev18_inR6 = {zll_main_dev84_in[2:0], zll_main_dev84_in[21:14], zll_main_dev84_in[13:11], zll_main_dev84_in[10:3], 3'h6};
  ZLL_Main_dev18  instR6 (zll_main_dev18_inR6[24:22], zll_main_dev18_inR6[21:14], zll_main_dev18_inR6[13:11], zll_main_dev18_inR6[10:3], zll_main_dev18_inR6[2:0], zll_main_dev18_outR6);
  assign zll_main_dev18_inR7 = {zll_main_dev84_in[2:0], zll_main_dev84_in[21:14], zll_main_dev84_in[13:11], zll_main_dev84_in[10:3], 3'h7};
  ZLL_Main_dev18  instR7 (zll_main_dev18_inR7[24:22], zll_main_dev18_inR7[21:14], zll_main_dev18_inR7[13:11], zll_main_dev18_inR7[10:3], zll_main_dev18_inR7[2:0], zll_main_dev18_outR7);
  assign zll_main_dev250_in = {zll_main_dev136_in[15:8], zll_main_dev136_in[7:0]};
  assign zll_main_dev253_in = {zll_main_dev250_in[15:8], zll_main_dev250_in[7:0]};
  assign zll_main_dev17_in = zll_main_dev253_in[15:0];
  assign zll_main_dev197_in = {zll_main_dev17_in[7:0], zll_main_dev17_in[15:8]};
  assign zll_main_dev3_in = {zll_main_dev197_in[15:8], zll_main_dev197_in[7:0], 3'h1};
  assign zll_main_dev69_in = {zll_main_dev3_in[18:11], zll_main_dev3_in[10:3], zll_main_dev3_in[2:0], 3'h2};
  assign zll_main_dev262_in = {3'h7, zll_main_dev69_in[2:0]};
  ZLL_Main_dev262  instR8 (zll_main_dev262_in[5:3], zll_main_dev262_in[2:0], zll_main_dev262_out);
  assign zll_main_dev252_in = {zll_main_dev69_in[21:14], zll_main_dev69_in[13:6], zll_main_dev69_in[5:3], zll_main_dev69_in[2:0], zll_main_dev262_out};
  assign zll_main_dev87_in = {zll_main_dev252_in[2:0], zll_main_dev252_in[16:9], zll_main_dev252_in[8:6], 1'h0};
  assign zll_main_dev176_in = {zll_main_dev87_in[14:12], zll_main_dev87_in[3:1], 1'h0};
  ZLL_Main_dev176  instR9 (zll_main_dev176_in[6:4], zll_main_dev176_in[3:1], zll_main_dev176_in[0], zll_main_dev176_out);
  assign id_in = {zll_main_dev87_in[14:12], zll_main_dev87_in[0]};
  assign zll_main_dev5_in = {zll_main_dev252_in[24:17], zll_main_dev252_in[16:9], zll_main_dev252_in[8:6], zll_main_dev252_in[5:3], (id_in[0] == 1'h1) ? id_in[3:1] : zll_main_dev176_out};
  assign zll_main_dev221_in = {zll_main_dev5_in[24:17], zll_main_dev5_in[16:9], zll_main_dev5_in[8:6], zll_main_dev5_in[5:3], zll_main_dev5_in[2:0], 3'h0};
  ZLL_Main_dev221  instR10 (zll_main_dev221_in[27:20], zll_main_dev221_in[19:12], zll_main_dev221_in[11:9], zll_main_dev221_in[8:6], zll_main_dev221_in[5:3], zll_main_dev221_in[2:0], zll_main_dev221_out);
  assign zll_main_dev221_inR1 = {zll_main_dev5_in[24:17], zll_main_dev5_in[16:9], zll_main_dev5_in[8:6], zll_main_dev5_in[5:3], zll_main_dev5_in[2:0], 3'h1};
  ZLL_Main_dev221  instR11 (zll_main_dev221_inR1[27:20], zll_main_dev221_inR1[19:12], zll_main_dev221_inR1[11:9], zll_main_dev221_inR1[8:6], zll_main_dev221_inR1[5:3], zll_main_dev221_inR1[2:0], zll_main_dev221_outR1);
  assign zll_main_dev221_inR2 = {zll_main_dev5_in[24:17], zll_main_dev5_in[16:9], zll_main_dev5_in[8:6], zll_main_dev5_in[5:3], zll_main_dev5_in[2:0], 3'h2};
  ZLL_Main_dev221  instR12 (zll_main_dev221_inR2[27:20], zll_main_dev221_inR2[19:12], zll_main_dev221_inR2[11:9], zll_main_dev221_inR2[8:6], zll_main_dev221_inR2[5:3], zll_main_dev221_inR2[2:0], zll_main_dev221_outR2);
  assign zll_main_dev221_inR3 = {zll_main_dev5_in[24:17], zll_main_dev5_in[16:9], zll_main_dev5_in[8:6], zll_main_dev5_in[5:3], zll_main_dev5_in[2:0], 3'h3};
  ZLL_Main_dev221  instR13 (zll_main_dev221_inR3[27:20], zll_main_dev221_inR3[19:12], zll_main_dev221_inR3[11:9], zll_main_dev221_inR3[8:6], zll_main_dev221_inR3[5:3], zll_main_dev221_inR3[2:0], zll_main_dev221_outR3);
  assign zll_main_dev221_inR4 = {zll_main_dev5_in[24:17], zll_main_dev5_in[16:9], zll_main_dev5_in[8:6], zll_main_dev5_in[5:3], zll_main_dev5_in[2:0], 3'h4};
  ZLL_Main_dev221  instR14 (zll_main_dev221_inR4[27:20], zll_main_dev221_inR4[19:12], zll_main_dev221_inR4[11:9], zll_main_dev221_inR4[8:6], zll_main_dev221_inR4[5:3], zll_main_dev221_inR4[2:0], zll_main_dev221_outR4);
  assign zll_main_dev221_inR5 = {zll_main_dev5_in[24:17], zll_main_dev5_in[16:9], zll_main_dev5_in[8:6], zll_main_dev5_in[5:3], zll_main_dev5_in[2:0], 3'h5};
  ZLL_Main_dev221  instR15 (zll_main_dev221_inR5[27:20], zll_main_dev221_inR5[19:12], zll_main_dev221_inR5[11:9], zll_main_dev221_inR5[8:6], zll_main_dev221_inR5[5:3], zll_main_dev221_inR5[2:0], zll_main_dev221_outR5);
  assign zll_main_dev221_inR6 = {zll_main_dev5_in[24:17], zll_main_dev5_in[16:9], zll_main_dev5_in[8:6], zll_main_dev5_in[5:3], zll_main_dev5_in[2:0], 3'h6};
  ZLL_Main_dev221  instR16 (zll_main_dev221_inR6[27:20], zll_main_dev221_inR6[19:12], zll_main_dev221_inR6[11:9], zll_main_dev221_inR6[8:6], zll_main_dev221_inR6[5:3], zll_main_dev221_inR6[2:0], zll_main_dev221_outR6);
  assign zll_main_dev221_inR7 = {zll_main_dev5_in[24:17], zll_main_dev5_in[16:9], zll_main_dev5_in[8:6], zll_main_dev5_in[5:3], zll_main_dev5_in[2:0], 3'h7};
  ZLL_Main_dev221  instR17 (zll_main_dev221_inR7[27:20], zll_main_dev221_inR7[19:12], zll_main_dev221_inR7[11:9], zll_main_dev221_inR7[8:6], zll_main_dev221_inR7[5:3], zll_main_dev221_inR7[2:0], zll_main_dev221_outR7);
  assign zll_main_dev142_in = {zll_main_dev136_in[15:8], zll_main_dev136_in[7:0]};
  assign zll_main_dev245_in = {zll_main_dev142_in[15:8], zll_main_dev142_in[7:0]};
  assign zll_main_dev99_in = zll_main_dev245_in[15:0];
  assign zll_main_dev120_in = {zll_main_dev99_in[7:0], zll_main_dev99_in[15:8]};
  assign zll_main_dev74_in = {zll_main_dev120_in[15:8], zll_main_dev120_in[7:0], 3'h1};
  assign zll_main_dev215_in = {zll_main_dev74_in[2:0], zll_main_dev74_in[18:11], zll_main_dev74_in[10:3]};
  assign zll_main_dev218_in = {zll_main_dev215_in[18:16], zll_main_dev215_in[15:8], zll_main_dev215_in[7:0], 3'h2};
  assign zll_main_dev262_inR1 = {3'h7, zll_main_dev218_in[2:0]};
  ZLL_Main_dev262  instR18 (zll_main_dev262_inR1[5:3], zll_main_dev262_inR1[2:0], zll_main_dev262_outR1);
  assign zll_main_dev125_in = {zll_main_dev218_in[21:19], zll_main_dev218_in[18:11], zll_main_dev218_in[2:0], zll_main_dev218_in[10:3], zll_main_dev262_outR1};
  assign zll_main_dev205_in = {zll_main_dev125_in[24:22], zll_main_dev125_in[2:0], zll_main_dev125_in[10:3], 1'h0};
  assign zll_main_dev103_in = {zll_main_dev205_in[14:12], zll_main_dev205_in[11:9], 1'h0};
  assign zll_main_dev285_in = {zll_main_dev103_in[6:4], zll_main_dev103_in[3:1], zll_main_dev103_in[0]};
  assign zll_main_dev270_in = {zll_main_dev285_in[3:1], zll_main_dev285_in[6:4]};
  ZLL_Main_dev270  instR19 (zll_main_dev270_in[5:3], zll_main_dev270_in[2:0], zll_main_dev270_out);
  assign id_inR1 = {zll_main_dev205_in[11:9], zll_main_dev205_in[0]};
  assign zll_main_dev202_in = {zll_main_dev125_in[21:14], zll_main_dev125_in[13:11], zll_main_dev125_in[10:3], (id_inR1[0] == 1'h1) ? id_inR1[3:1] : zll_main_dev270_out};
  assign zll_main_dev101_in = {zll_main_dev202_in[21:14], zll_main_dev202_in[13:11], zll_main_dev202_in[2:0], zll_main_dev202_in[10:3], 3'h0};
  ZLL_Main_dev101  instR20 (zll_main_dev101_in[24:17], zll_main_dev101_in[16:14], zll_main_dev101_in[13:11], zll_main_dev101_in[10:3], zll_main_dev101_in[2:0], zll_main_dev101_out);
  assign zll_main_dev101_inR1 = {zll_main_dev202_in[21:14], zll_main_dev202_in[13:11], zll_main_dev202_in[2:0], zll_main_dev202_in[10:3], 3'h1};
  ZLL_Main_dev101  instR21 (zll_main_dev101_inR1[24:17], zll_main_dev101_inR1[16:14], zll_main_dev101_inR1[13:11], zll_main_dev101_inR1[10:3], zll_main_dev101_inR1[2:0], zll_main_dev101_outR1);
  assign zll_main_dev101_inR2 = {zll_main_dev202_in[21:14], zll_main_dev202_in[13:11], zll_main_dev202_in[2:0], zll_main_dev202_in[10:3], 3'h2};
  ZLL_Main_dev101  instR22 (zll_main_dev101_inR2[24:17], zll_main_dev101_inR2[16:14], zll_main_dev101_inR2[13:11], zll_main_dev101_inR2[10:3], zll_main_dev101_inR2[2:0], zll_main_dev101_outR2);
  assign zll_main_dev101_inR3 = {zll_main_dev202_in[21:14], zll_main_dev202_in[13:11], zll_main_dev202_in[2:0], zll_main_dev202_in[10:3], 3'h3};
  ZLL_Main_dev101  instR23 (zll_main_dev101_inR3[24:17], zll_main_dev101_inR3[16:14], zll_main_dev101_inR3[13:11], zll_main_dev101_inR3[10:3], zll_main_dev101_inR3[2:0], zll_main_dev101_outR3);
  assign zll_main_dev101_inR4 = {zll_main_dev202_in[21:14], zll_main_dev202_in[13:11], zll_main_dev202_in[2:0], zll_main_dev202_in[10:3], 3'h4};
  ZLL_Main_dev101  instR24 (zll_main_dev101_inR4[24:17], zll_main_dev101_inR4[16:14], zll_main_dev101_inR4[13:11], zll_main_dev101_inR4[10:3], zll_main_dev101_inR4[2:0], zll_main_dev101_outR4);
  assign zll_main_dev101_inR5 = {zll_main_dev202_in[21:14], zll_main_dev202_in[13:11], zll_main_dev202_in[2:0], zll_main_dev202_in[10:3], 3'h5};
  ZLL_Main_dev101  instR25 (zll_main_dev101_inR5[24:17], zll_main_dev101_inR5[16:14], zll_main_dev101_inR5[13:11], zll_main_dev101_inR5[10:3], zll_main_dev101_inR5[2:0], zll_main_dev101_outR5);
  assign zll_main_dev101_inR6 = {zll_main_dev202_in[21:14], zll_main_dev202_in[13:11], zll_main_dev202_in[2:0], zll_main_dev202_in[10:3], 3'h6};
  ZLL_Main_dev101  instR26 (zll_main_dev101_inR6[24:17], zll_main_dev101_inR6[16:14], zll_main_dev101_inR6[13:11], zll_main_dev101_inR6[10:3], zll_main_dev101_inR6[2:0], zll_main_dev101_outR6);
  assign zll_main_dev101_inR7 = {zll_main_dev202_in[21:14], zll_main_dev202_in[13:11], zll_main_dev202_in[2:0], zll_main_dev202_in[10:3], 3'h7};
  ZLL_Main_dev101  instR27 (zll_main_dev101_inR7[24:17], zll_main_dev101_inR7[16:14], zll_main_dev101_inR7[13:11], zll_main_dev101_inR7[10:3], zll_main_dev101_inR7[2:0], zll_main_dev101_outR7);
  assign zll_main_dev234_in = {zll_main_dev136_in[15:8], zll_main_dev136_in[7:0]};
  assign zll_main_dev38_in = {zll_main_dev234_in[15:8], zll_main_dev234_in[7:0]};
  assign zll_main_dev169_in = zll_main_dev38_in[15:0];
  assign zll_main_dev37_in = {zll_main_dev169_in[15:8], zll_main_dev169_in[7:0], 3'h1};
  assign zll_main_dev42_in = {zll_main_dev37_in[18:11], zll_main_dev37_in[10:3], zll_main_dev37_in[2:0], 3'h2};
  assign zll_main_dev262_inR2 = {3'h7, zll_main_dev42_in[2:0]};
  ZLL_Main_dev262  instR28 (zll_main_dev262_inR2[5:3], zll_main_dev262_inR2[2:0], zll_main_dev262_outR2);
  assign zll_main_dev171_in = {zll_main_dev42_in[21:14], zll_main_dev42_in[2:0], zll_main_dev42_in[13:6], zll_main_dev42_in[5:3], zll_main_dev262_outR2};
  assign zll_main_dev89_in = {zll_main_dev171_in[24:17], zll_main_dev171_in[2:0], zll_main_dev171_in[5:3], 1'h0};
  assign zll_main_dev176_inR1 = {zll_main_dev89_in[6:4], zll_main_dev89_in[3:1], 1'h0};
  ZLL_Main_dev176  instR29 (zll_main_dev176_inR1[6:4], zll_main_dev176_inR1[3:1], zll_main_dev176_inR1[0], zll_main_dev176_outR1);
  assign id_inR2 = {zll_main_dev89_in[6:4], zll_main_dev89_in[0]};
  assign zll_main_dev27_in = {zll_main_dev171_in[24:17], zll_main_dev171_in[16:14], zll_main_dev171_in[13:6], zll_main_dev171_in[5:3], (id_inR2[0] == 1'h1) ? id_inR2[3:1] : zll_main_dev176_outR1};
  assign zll_main_dev272_in = {zll_main_dev27_in[24:17], zll_main_dev27_in[16:14], zll_main_dev27_in[13:6], zll_main_dev27_in[5:3], zll_main_dev27_in[2:0], 3'h0};
  ZLL_Main_dev272  instR30 (zll_main_dev272_in[27:20], zll_main_dev272_in[19:17], zll_main_dev272_in[16:9], zll_main_dev272_in[8:6], zll_main_dev272_in[5:3], zll_main_dev272_in[2:0], zll_main_dev272_out);
  assign zll_main_dev272_inR1 = {zll_main_dev27_in[24:17], zll_main_dev27_in[16:14], zll_main_dev27_in[13:6], zll_main_dev27_in[5:3], zll_main_dev27_in[2:0], 3'h1};
  ZLL_Main_dev272  instR31 (zll_main_dev272_inR1[27:20], zll_main_dev272_inR1[19:17], zll_main_dev272_inR1[16:9], zll_main_dev272_inR1[8:6], zll_main_dev272_inR1[5:3], zll_main_dev272_inR1[2:0], zll_main_dev272_outR1);
  assign zll_main_dev272_inR2 = {zll_main_dev27_in[24:17], zll_main_dev27_in[16:14], zll_main_dev27_in[13:6], zll_main_dev27_in[5:3], zll_main_dev27_in[2:0], 3'h2};
  ZLL_Main_dev272  instR32 (zll_main_dev272_inR2[27:20], zll_main_dev272_inR2[19:17], zll_main_dev272_inR2[16:9], zll_main_dev272_inR2[8:6], zll_main_dev272_inR2[5:3], zll_main_dev272_inR2[2:0], zll_main_dev272_outR2);
  assign zll_main_dev272_inR3 = {zll_main_dev27_in[24:17], zll_main_dev27_in[16:14], zll_main_dev27_in[13:6], zll_main_dev27_in[5:3], zll_main_dev27_in[2:0], 3'h3};
  ZLL_Main_dev272  instR33 (zll_main_dev272_inR3[27:20], zll_main_dev272_inR3[19:17], zll_main_dev272_inR3[16:9], zll_main_dev272_inR3[8:6], zll_main_dev272_inR3[5:3], zll_main_dev272_inR3[2:0], zll_main_dev272_outR3);
  assign zll_main_dev272_inR4 = {zll_main_dev27_in[24:17], zll_main_dev27_in[16:14], zll_main_dev27_in[13:6], zll_main_dev27_in[5:3], zll_main_dev27_in[2:0], 3'h4};
  ZLL_Main_dev272  instR34 (zll_main_dev272_inR4[27:20], zll_main_dev272_inR4[19:17], zll_main_dev272_inR4[16:9], zll_main_dev272_inR4[8:6], zll_main_dev272_inR4[5:3], zll_main_dev272_inR4[2:0], zll_main_dev272_outR4);
  assign zll_main_dev272_inR5 = {zll_main_dev27_in[24:17], zll_main_dev27_in[16:14], zll_main_dev27_in[13:6], zll_main_dev27_in[5:3], zll_main_dev27_in[2:0], 3'h5};
  ZLL_Main_dev272  instR35 (zll_main_dev272_inR5[27:20], zll_main_dev272_inR5[19:17], zll_main_dev272_inR5[16:9], zll_main_dev272_inR5[8:6], zll_main_dev272_inR5[5:3], zll_main_dev272_inR5[2:0], zll_main_dev272_outR5);
  assign zll_main_dev272_inR6 = {zll_main_dev27_in[24:17], zll_main_dev27_in[16:14], zll_main_dev27_in[13:6], zll_main_dev27_in[5:3], zll_main_dev27_in[2:0], 3'h6};
  ZLL_Main_dev272  instR36 (zll_main_dev272_inR6[27:20], zll_main_dev272_inR6[19:17], zll_main_dev272_inR6[16:9], zll_main_dev272_inR6[8:6], zll_main_dev272_inR6[5:3], zll_main_dev272_inR6[2:0], zll_main_dev272_outR6);
  assign zll_main_dev272_inR7 = {zll_main_dev27_in[24:17], zll_main_dev27_in[16:14], zll_main_dev27_in[13:6], zll_main_dev27_in[5:3], zll_main_dev27_in[2:0], 3'h7};
  ZLL_Main_dev272  instR37 (zll_main_dev272_inR7[27:20], zll_main_dev272_inR7[19:17], zll_main_dev272_inR7[16:9], zll_main_dev272_inR7[8:6], zll_main_dev272_inR7[5:3], zll_main_dev272_inR7[2:0], zll_main_dev272_outR7);
  assign {__continue, __out0, __out1, __out2, __out3} = {{zll_main_dev18_out, zll_main_dev18_outR1, zll_main_dev18_outR2, zll_main_dev18_outR3, zll_main_dev18_outR4, zll_main_dev18_outR5, zll_main_dev18_outR6, zll_main_dev18_outR7}, {zll_main_dev221_out, zll_main_dev221_outR1, zll_main_dev221_outR2, zll_main_dev221_outR3, zll_main_dev221_outR4, zll_main_dev221_outR5, zll_main_dev221_outR6, zll_main_dev221_outR7}, {zll_main_dev101_out, zll_main_dev101_outR1, zll_main_dev101_outR2, zll_main_dev101_outR3, zll_main_dev101_outR4, zll_main_dev101_outR5, zll_main_dev101_outR6, zll_main_dev101_outR7}, {zll_main_dev272_out, zll_main_dev272_outR1, zll_main_dev272_outR2, zll_main_dev272_outR3, zll_main_dev272_outR4, zll_main_dev272_outR5, zll_main_dev272_outR6, zll_main_dev272_outR7}};
endmodule

module ZLL_Main_dev280 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  output logic [2:0] res);
  logic [5:0] zll_main_dev282_in;
  logic [5:0] zll_main_dev159_in;
  logic [2:0] resize_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR2;
  assign zll_main_dev282_in = {arg0, arg1};
  assign zll_main_dev159_in = zll_main_dev282_in[5:0];
  assign resize_in = zll_main_dev159_in[5:3];
  assign resize_inR1 = zll_main_dev159_in[2:0];
  assign binop_in = {128'(resize_in[2:0]), 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h8};
  assign resize_inR2 = binop_inR1[255:128] % binop_inR1[127:0];
  assign res = resize_inR2[2:0];
endmodule

module ZLL_Main_dev272 (input logic [7:0] arg0,
  input logic [2:0] arg1,
  input logic [7:0] arg2,
  input logic [2:0] arg3,
  input logic [2:0] arg4,
  input logic [2:0] arg5,
  output logic [0:0] res);
  logic [5:0] zll_main_dev198_in;
  logic [0:0] zll_main_dev198_out;
  logic [28:0] zll_main_dev124_in;
  logic [5:0] zll_main_dev198_inR1;
  logic [0:0] zll_main_dev198_outR1;
  logic [20:0] zll_main_dev93_in;
  logic [20:0] zll_main_dev199_in;
  logic [7:0] resize_in;
  logic [5:0] zll_main_dev280_in;
  logic [2:0] zll_main_dev280_out;
  logic [5:0] zll_main_dev214_in;
  logic [2:0] zll_main_dev214_out;
  logic [5:0] zll_main_dev270_in;
  logic [2:0] zll_main_dev270_out;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR2;
  logic [17:0] zll_main_dev102_in;
  logic [7:0] resize_inR3;
  logic [5:0] zll_main_dev214_inR1;
  logic [2:0] zll_main_dev214_outR1;
  logic [5:0] zll_main_dev270_inR1;
  logic [2:0] zll_main_dev270_outR1;
  logic [2:0] resize_inR4;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR5;
  assign zll_main_dev198_in = {arg5, arg4};
  ZLL_Main_dev198  inst (zll_main_dev198_in[5:3], zll_main_dev198_in[2:0], zll_main_dev198_out);
  assign zll_main_dev124_in = {arg0, arg1, arg2, arg3, arg5, arg4, zll_main_dev198_out};
  assign zll_main_dev198_inR1 = {zll_main_dev124_in[6:4], zll_main_dev124_in[3:1]};
  ZLL_Main_dev198  instR1 (zll_main_dev198_inR1[5:3], zll_main_dev198_inR1[2:0], zll_main_dev198_outR1);
  assign zll_main_dev93_in = {zll_main_dev124_in[20:18], zll_main_dev124_in[17:10], zll_main_dev124_in[9:7], zll_main_dev124_in[6:4], zll_main_dev124_in[3:1], zll_main_dev198_outR1};
  assign zll_main_dev199_in = {zll_main_dev93_in[20:18], zll_main_dev93_in[17:10], zll_main_dev93_in[9:7], zll_main_dev93_in[6:4], zll_main_dev93_in[3:1], zll_main_dev93_in[0]};
  assign resize_in = zll_main_dev199_in[17:10];
  assign zll_main_dev280_in = {zll_main_dev199_in[6:4], zll_main_dev199_in[3:1]};
  ZLL_Main_dev280  instR2 (zll_main_dev280_in[5:3], zll_main_dev280_in[2:0], zll_main_dev280_out);
  assign zll_main_dev214_in = {zll_main_dev280_out, zll_main_dev199_in[20:18]};
  ZLL_Main_dev214  instR3 (zll_main_dev214_in[5:3], zll_main_dev214_in[2:0], zll_main_dev214_out);
  assign zll_main_dev270_in = {zll_main_dev214_out, zll_main_dev199_in[9:7]};
  ZLL_Main_dev270  instR4 (zll_main_dev270_in[5:3], zll_main_dev270_in[2:0], zll_main_dev270_out);
  assign resize_inR1 = zll_main_dev270_out;
  assign binop_in = {128'h8, 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h1};
  assign binop_inR3 = {128'(resize_in[7:0]), binop_inR2[255:128] * binop_inR2[127:0]};
  assign resize_inR2 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign zll_main_dev102_in = {zll_main_dev124_in[28:21], zll_main_dev124_in[20:18], zll_main_dev124_in[9:7], zll_main_dev124_in[6:4], zll_main_dev124_in[0]};
  assign resize_inR3 = zll_main_dev102_in[17:10];
  assign zll_main_dev214_inR1 = {zll_main_dev102_in[3:1], zll_main_dev102_in[9:7]};
  ZLL_Main_dev214  instR5 (zll_main_dev214_inR1[5:3], zll_main_dev214_inR1[2:0], zll_main_dev214_outR1);
  assign zll_main_dev270_inR1 = {zll_main_dev214_outR1, zll_main_dev102_in[6:4]};
  ZLL_Main_dev270  instR6 (zll_main_dev270_inR1[5:3], zll_main_dev270_inR1[2:0], zll_main_dev270_outR1);
  assign resize_inR4 = zll_main_dev270_outR1;
  assign binop_inR4 = {128'h8, 128'(resize_inR4[2:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h1};
  assign binop_inR7 = {128'(resize_inR3[7:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR5 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign res = (zll_main_dev102_in[0] == 1'h1) ? resize_inR5[0] : resize_inR2[0];
endmodule

module ZLL_Main_dev270 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  output logic [2:0] res);
  logic [5:0] zll_main_dev228_in;
  logic [5:0] zll_main_dev276_in;
  logic [2:0] resize_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR2;
  assign zll_main_dev228_in = {arg0, arg1};
  assign zll_main_dev276_in = zll_main_dev228_in[5:0];
  assign resize_in = zll_main_dev276_in[5:3];
  assign resize_inR1 = zll_main_dev276_in[2:0];
  assign binop_in = {128'(resize_in[2:0]), 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] + binop_in[127:0], 128'h8};
  assign resize_inR2 = binop_inR1[255:128] % binop_inR1[127:0];
  assign res = resize_inR2[2:0];
endmodule

module ZLL_Main_dev262 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  output logic [2:0] res);
  logic [5:0] zll_main_dev208_in;
  logic [5:0] zll_main_dev258_in;
  logic [2:0] resize_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR2;
  assign zll_main_dev208_in = {arg0, arg1};
  assign zll_main_dev258_in = zll_main_dev208_in[5:0];
  assign resize_in = zll_main_dev258_in[5:3];
  assign resize_inR1 = zll_main_dev258_in[2:0];
  assign binop_in = {128'(resize_in[2:0]), 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] / binop_in[127:0], 128'h8};
  assign resize_inR2 = binop_inR1[255:128] % binop_inR1[127:0];
  assign res = resize_inR2[2:0];
endmodule

module ZLL_Main_dev229 (input logic [2:0] arg0,
  output logic [0:0] res);
  logic [2:0] resize_in;
  logic [127:0] zll_main_dev187_in;
  logic [127:0] resize_inR1;
  logic [0:0] msbit_in;
  logic [0:0] rewire_prelude_not_in;
  logic [1:0] zll_rewire_prelude_not_in;
  logic [0:0] lit_in;
  assign resize_in = arg0;
  assign zll_main_dev187_in = 128'(resize_in[2:0]);
  assign resize_inR1 = zll_main_dev187_in[127:0];
  assign msbit_in = resize_inR1[0];
  assign rewire_prelude_not_in = msbit_in[0];
  assign zll_rewire_prelude_not_in = {rewire_prelude_not_in[0], rewire_prelude_not_in[0]};
  assign lit_in = zll_rewire_prelude_not_in[0];
  assign res = (lit_in[0] == 1'h1) ? 1'h0 : 1'h1;
endmodule

module ZLL_Main_dev221 (input logic [7:0] arg0,
  input logic [7:0] arg1,
  input logic [2:0] arg2,
  input logic [2:0] arg3,
  input logic [2:0] arg4,
  input logic [2:0] arg5,
  output logic [0:0] res);
  logic [2:0] zll_main_dev229_in;
  logic [0:0] zll_main_dev229_out;
  logic [28:0] zll_main_dev122_in;
  logic [2:0] zll_main_dev229_inR1;
  logic [0:0] zll_main_dev229_outR1;
  logic [20:0] zll_main_dev81_in;
  logic [20:0] zll_main_dev150_in;
  logic [7:0] resize_in;
  logic [5:0] zll_main_dev280_in;
  logic [2:0] zll_main_dev280_out;
  logic [5:0] zll_main_dev262_in;
  logic [2:0] zll_main_dev262_out;
  logic [5:0] zll_main_dev270_in;
  logic [2:0] zll_main_dev270_out;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR2;
  logic [17:0] zll_main_dev235_in;
  logic [7:0] resize_inR3;
  logic [5:0] zll_main_dev262_inR1;
  logic [2:0] zll_main_dev262_outR1;
  logic [5:0] zll_main_dev270_inR1;
  logic [2:0] zll_main_dev270_outR1;
  logic [2:0] resize_inR4;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR5;
  assign zll_main_dev229_in = arg5;
  ZLL_Main_dev229  inst (zll_main_dev229_in[2:0], zll_main_dev229_out);
  assign zll_main_dev122_in = {arg0, arg5, arg1, arg2, arg3, arg4, zll_main_dev229_out};
  assign zll_main_dev229_inR1 = zll_main_dev122_in[20:18];
  ZLL_Main_dev229  instR1 (zll_main_dev229_inR1[2:0], zll_main_dev229_outR1);
  assign zll_main_dev81_in = {zll_main_dev122_in[28:21], zll_main_dev122_in[20:18], zll_main_dev122_in[9:7], zll_main_dev122_in[6:4], zll_main_dev122_in[3:1], zll_main_dev229_outR1};
  assign zll_main_dev150_in = {zll_main_dev81_in[20:13], zll_main_dev81_in[12:10], zll_main_dev81_in[9:7], zll_main_dev81_in[6:4], zll_main_dev81_in[3:1], zll_main_dev81_in[0]};
  assign resize_in = zll_main_dev150_in[20:13];
  assign zll_main_dev280_in = {zll_main_dev150_in[12:10], zll_main_dev150_in[9:7]};
  ZLL_Main_dev280  instR2 (zll_main_dev280_in[5:3], zll_main_dev280_in[2:0], zll_main_dev280_out);
  assign zll_main_dev262_in = {zll_main_dev280_out, zll_main_dev150_in[6:4]};
  ZLL_Main_dev262  instR3 (zll_main_dev262_in[5:3], zll_main_dev262_in[2:0], zll_main_dev262_out);
  assign zll_main_dev270_in = {zll_main_dev150_in[3:1], zll_main_dev262_out};
  ZLL_Main_dev270  instR4 (zll_main_dev270_in[5:3], zll_main_dev270_in[2:0], zll_main_dev270_out);
  assign resize_inR1 = zll_main_dev270_out;
  assign binop_in = {128'h8, 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h1};
  assign binop_inR3 = {128'(resize_in[7:0]), binop_inR2[255:128] * binop_inR2[127:0]};
  assign resize_inR2 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign zll_main_dev235_in = {zll_main_dev122_in[20:18], zll_main_dev122_in[17:10], zll_main_dev122_in[6:4], zll_main_dev122_in[3:1], zll_main_dev122_in[0]};
  assign resize_inR3 = zll_main_dev235_in[14:7];
  assign zll_main_dev262_inR1 = {zll_main_dev235_in[17:15], zll_main_dev235_in[6:4]};
  ZLL_Main_dev262  instR5 (zll_main_dev262_inR1[5:3], zll_main_dev262_inR1[2:0], zll_main_dev262_outR1);
  assign zll_main_dev270_inR1 = {zll_main_dev235_in[3:1], zll_main_dev262_outR1};
  ZLL_Main_dev270  instR6 (zll_main_dev270_inR1[5:3], zll_main_dev270_inR1[2:0], zll_main_dev270_outR1);
  assign resize_inR4 = zll_main_dev270_outR1;
  assign binop_inR4 = {128'h8, 128'(resize_inR4[2:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h1};
  assign binop_inR7 = {128'(resize_inR3[7:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR5 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign res = (zll_main_dev235_in[0] == 1'h1) ? resize_inR5[0] : resize_inR2[0];
endmodule

module ZLL_Main_dev214 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  output logic [2:0] res);
  logic [5:0] zll_main_dev274_in;
  logic [5:0] zll_main_dev112_in;
  logic [2:0] resize_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR2;
  assign zll_main_dev274_in = {arg0, arg1};
  assign zll_main_dev112_in = zll_main_dev274_in[5:0];
  assign resize_in = zll_main_dev112_in[5:3];
  assign resize_inR1 = zll_main_dev112_in[2:0];
  assign binop_in = {128'(resize_in[2:0]), 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] * binop_in[127:0], 128'h8};
  assign resize_inR2 = binop_inR1[255:128] % binop_inR1[127:0];
  assign res = resize_inR2[2:0];
endmodule

module ZLL_Main_dev198 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  output logic [0:0] res);
  logic [5:0] zll_main_dev145_in;
  logic [5:0] zll_main_dev217_in;
  logic [2:0] resize_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  assign zll_main_dev145_in = {arg0, arg1};
  assign zll_main_dev217_in = zll_main_dev145_in[5:0];
  assign resize_in = zll_main_dev217_in[5:3];
  assign resize_inR1 = zll_main_dev217_in[2:0];
  assign binop_in = {128'(resize_in[2:0]), 128'(resize_inR1[2:0])};
  assign res = binop_in[255:128] < binop_in[127:0];
endmodule

module ZLL_Main_dev176 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  input logic [0:0] arg2,
  output logic [2:0] res);
  logic [6:0] zll_main_dev211_in;
  logic [5:0] zll_main_dev270_in;
  logic [2:0] zll_main_dev270_out;
  assign zll_main_dev211_in = {arg0, arg1, arg2};
  assign zll_main_dev270_in = {zll_main_dev211_in[6:4], zll_main_dev211_in[3:1]};
  ZLL_Main_dev270  inst (zll_main_dev270_in[5:3], zll_main_dev270_in[2:0], zll_main_dev270_out);
  assign res = zll_main_dev270_out;
endmodule

module ZLL_Main_dev101 (input logic [7:0] arg0,
  input logic [2:0] arg1,
  input logic [2:0] arg2,
  input logic [7:0] arg3,
  input logic [2:0] arg4,
  output logic [0:0] res);
  logic [5:0] zll_main_dev198_in;
  logic [0:0] zll_main_dev198_out;
  logic [25:0] zll_main_dev107_in;
  logic [5:0] zll_main_dev198_inR1;
  logic [0:0] zll_main_dev198_outR1;
  logic [17:0] zll_main_dev267_in;
  logic [17:0] zll_main_dev219_in;
  logic [7:0] resize_in;
  logic [5:0] zll_main_dev280_in;
  logic [2:0] zll_main_dev280_out;
  logic [5:0] zll_main_dev214_in;
  logic [2:0] zll_main_dev214_out;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR2;
  logic [14:0] zll_main_dev131_in;
  logic [7:0] resize_inR3;
  logic [5:0] zll_main_dev214_inR1;
  logic [2:0] zll_main_dev214_outR1;
  logic [2:0] resize_inR4;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR5;
  assign zll_main_dev198_in = {arg4, arg2};
  ZLL_Main_dev198  inst (zll_main_dev198_in[5:3], zll_main_dev198_in[2:0], zll_main_dev198_out);
  assign zll_main_dev107_in = {arg0, arg1, arg2, arg4, arg3, zll_main_dev198_out};
  assign zll_main_dev198_inR1 = {zll_main_dev107_in[11:9], zll_main_dev107_in[14:12]};
  ZLL_Main_dev198  instR1 (zll_main_dev198_inR1[5:3], zll_main_dev198_inR1[2:0], zll_main_dev198_outR1);
  assign zll_main_dev267_in = {zll_main_dev107_in[25:18], zll_main_dev107_in[17:15], zll_main_dev107_in[14:12], zll_main_dev107_in[11:9], zll_main_dev198_outR1};
  assign zll_main_dev219_in = {zll_main_dev267_in[17:10], zll_main_dev267_in[9:7], zll_main_dev267_in[6:4], zll_main_dev267_in[3:1], zll_main_dev267_in[0]};
  assign resize_in = zll_main_dev219_in[17:10];
  assign zll_main_dev280_in = {zll_main_dev219_in[3:1], zll_main_dev219_in[6:4]};
  ZLL_Main_dev280  instR2 (zll_main_dev280_in[5:3], zll_main_dev280_in[2:0], zll_main_dev280_out);
  assign zll_main_dev214_in = {zll_main_dev280_out, zll_main_dev219_in[9:7]};
  ZLL_Main_dev214  instR3 (zll_main_dev214_in[5:3], zll_main_dev214_in[2:0], zll_main_dev214_out);
  assign resize_inR1 = zll_main_dev214_out;
  assign binop_in = {128'h8, 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h1};
  assign binop_inR3 = {128'(resize_in[7:0]), binop_inR2[255:128] * binop_inR2[127:0]};
  assign resize_inR2 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign zll_main_dev131_in = {zll_main_dev107_in[17:15], zll_main_dev107_in[11:9], zll_main_dev107_in[8:1], zll_main_dev107_in[0]};
  assign resize_inR3 = zll_main_dev131_in[8:1];
  assign zll_main_dev214_inR1 = {zll_main_dev131_in[11:9], zll_main_dev131_in[14:12]};
  ZLL_Main_dev214  instR4 (zll_main_dev214_inR1[5:3], zll_main_dev214_inR1[2:0], zll_main_dev214_outR1);
  assign resize_inR4 = zll_main_dev214_outR1;
  assign binop_inR4 = {128'h8, 128'(resize_inR4[2:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h1};
  assign binop_inR7 = {128'(resize_inR3[7:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR5 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign res = (zll_main_dev131_in[0] == 1'h1) ? resize_inR5[0] : resize_inR2[0];
endmodule

module ZLL_Main_dev18 (input logic [2:0] arg0,
  input logic [7:0] arg1,
  input logic [2:0] arg2,
  input logic [7:0] arg3,
  input logic [2:0] arg4,
  output logic [0:0] res);
  logic [2:0] zll_main_dev229_in;
  logic [0:0] zll_main_dev229_out;
  logic [25:0] zll_main_dev30_in;
  logic [2:0] zll_main_dev229_inR1;
  logic [0:0] zll_main_dev229_outR1;
  logic [17:0] zll_main_dev203_in;
  logic [17:0] zll_main_dev263_in;
  logic [7:0] resize_in;
  logic [5:0] zll_main_dev280_in;
  logic [2:0] zll_main_dev280_out;
  logic [5:0] zll_main_dev262_in;
  logic [2:0] zll_main_dev262_out;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR2;
  logic [14:0] zll_main_dev_in;
  logic [7:0] resize_inR3;
  logic [5:0] zll_main_dev262_inR1;
  logic [2:0] zll_main_dev262_outR1;
  logic [2:0] resize_inR4;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR5;
  assign zll_main_dev229_in = arg4;
  ZLL_Main_dev229  inst (zll_main_dev229_in[2:0], zll_main_dev229_out);
  assign zll_main_dev30_in = {arg4, arg0, arg1, arg2, arg3, zll_main_dev229_out};
  assign zll_main_dev229_inR1 = zll_main_dev30_in[25:23];
  ZLL_Main_dev229  instR1 (zll_main_dev229_inR1[2:0], zll_main_dev229_outR1);
  assign zll_main_dev203_in = {zll_main_dev30_in[25:23], zll_main_dev30_in[22:20], zll_main_dev30_in[11:9], zll_main_dev30_in[8:1], zll_main_dev229_outR1};
  assign zll_main_dev263_in = {zll_main_dev203_in[17:15], zll_main_dev203_in[14:12], zll_main_dev203_in[11:9], zll_main_dev203_in[8:1], zll_main_dev203_in[0]};
  assign resize_in = zll_main_dev263_in[8:1];
  assign zll_main_dev280_in = {zll_main_dev263_in[17:15], zll_main_dev263_in[11:9]};
  ZLL_Main_dev280  instR2 (zll_main_dev280_in[5:3], zll_main_dev280_in[2:0], zll_main_dev280_out);
  assign zll_main_dev262_in = {zll_main_dev280_out, zll_main_dev263_in[14:12]};
  ZLL_Main_dev262  instR3 (zll_main_dev262_in[5:3], zll_main_dev262_in[2:0], zll_main_dev262_out);
  assign resize_inR1 = zll_main_dev262_out;
  assign binop_in = {128'h8, 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h1};
  assign binop_inR3 = {128'(resize_in[7:0]), binop_inR2[255:128] * binop_inR2[127:0]};
  assign resize_inR2 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign zll_main_dev_in = {zll_main_dev30_in[25:23], zll_main_dev30_in[22:20], zll_main_dev30_in[19:12], zll_main_dev30_in[0]};
  assign resize_inR3 = zll_main_dev_in[8:1];
  assign zll_main_dev262_inR1 = {zll_main_dev_in[14:12], zll_main_dev_in[11:9]};
  ZLL_Main_dev262  instR4 (zll_main_dev262_inR1[5:3], zll_main_dev262_inR1[2:0], zll_main_dev262_outR1);
  assign resize_inR4 = zll_main_dev262_outR1;
  assign binop_inR4 = {128'h8, 128'(resize_inR4[2:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h1};
  assign binop_inR7 = {128'(resize_inR3[7:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR5 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign res = (zll_main_dev_in[0] == 1'h1) ? resize_inR5[0] : resize_inR2[0];
endmodule