module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [9:0] __in0,
  output logic [15:0] __out0);
  logic [39:0] rewire_monad_iterst_in;
  logic [69:0] zll_rewire_monad_iterst_in;
  logic [69:0] zll_rewire_monad_iterst32_in;
  logic [39:0] main_loop_in;
  logic [39:0] zll_main_loop3_in;
  logic [39:0] zll_main_loop6_in;
  logic [29:0] zll_main_loop5_in;
  logic [29:0] id_in;
  logic [24:0] main_inputtomystate_in;
  logic [49:0] zll_main_inputtomystate_in;
  logic [49:0] zll_main_inputtomystate18_in;
  logic [49:0] zll_main_inputtomystate17_in;
  logic [49:0] zll_main_inputtomystate9_in;
  logic [24:0] zll_main_inputtomystate1_in;
  logic [24:0] zll_main_inputtomystate3_in;
  logic [13:0] zll_main_inputtomystate12_in;
  logic [24:0] zll_main_inputtomystate14_in;
  logic [24:0] zll_main_inputtomystate13_in;
  logic [12:0] zll_main_inputtomystate8_in;
  logic [24:0] zll_main_inputtomystate16_in;
  logic [22:0] zll_main_inputtomystate2_in;
  logic [24:0] zll_main_inputtomystate10_in;
  logic [18:0] zll_main_inputtomystate11_in;
  logic [13:0] zll_main_inputtomystate15_in;
  logic [44:0] zll_main_incrpipeline5_in;
  logic [44:0] zll_main_incrpipeline4_in;
  logic [29:0] id_inR1;
  logic [29:0] zll_main_incrpipeline8_in;
  logic [29:0] zll_main_incrpipeline6_in;
  logic [29:0] id_inR2;
  logic [29:0] zll_main_incrpipeline10_in;
  logic [29:0] resize_in;
  logic [255:0] binop_in;
  logic [127:0] resize_inR1;
  logic [44:0] zll_main_loop1_in;
  logic [44:0] zll_main_loop4_in;
  logic [14:0] main_mystatetooutput_in;
  logic [29:0] zll_main_mystatetooutput4_in;
  logic [29:0] zll_main_mystatetooutput7_in;
  logic [14:0] zll_main_mystatetooutput1_in;
  logic [14:0] zll_main_mystatetooutput3_in;
  logic [8:0] zll_main_mystatetooutput_in;
  logic [14:0] zll_main_mystatetooutput2_in;
  logic [12:0] zll_main_mystatetooutput8_in;
  logic [14:0] zll_main_mystatetooutput5_in;
  logic [8:0] zll_main_mystatetooutput6_in;
  logic [75:0] zll_rewire_monad_iterst27_in;
  logic [75:0] zll_rewire_monad_iterst25_in;
  logic [77:0] zll_rewire_monad_iterst36_in;
  logic [77:0] zll_rewire_monad_iterst26_in;
  logic [75:0] zll_rewire_monad_iterst35_in;
  logic [75:0] zll_rewire_monad_iterst22_in;
  logic [75:0] zll_rewire_monad_iterst37_in;
  logic [75:0] zll_rewire_monad_iterst31_in;
  logic [29:0] zll_rewire_monad_iterst15_in;
  logic [93:0] zll_rewire_monad_iterst4_in;
  logic [93:0] zll_rewire_monad_iterst29_in;
  logic [45:0] zll_rewire_monad_iterst33_in;
  logic [31:0] __padding;
  logic [29:0] __st0;
  logic [29:0] __st0_next;
  assign rewire_monad_iterst_in = {__in0, __st0};
  assign zll_rewire_monad_iterst_in = {rewire_monad_iterst_in[39:30], rewire_monad_iterst_in[29:0], rewire_monad_iterst_in[29:0]};
  assign zll_rewire_monad_iterst32_in = {zll_rewire_monad_iterst_in[69:60], zll_rewire_monad_iterst_in[59:0]};
  assign main_loop_in = {zll_rewire_monad_iterst32_in[69:60], zll_rewire_monad_iterst32_in[59:30]};
  assign zll_main_loop3_in = {main_loop_in[39:30], main_loop_in[29:0]};
  assign zll_main_loop6_in = zll_main_loop3_in[39:0];
  assign zll_main_loop5_in = zll_main_loop6_in[29:0];
  assign id_in = zll_main_loop5_in[29:0];
  assign main_inputtomystate_in = {zll_main_loop6_in[39:30], id_in[29:15]};
  assign zll_main_inputtomystate_in = {main_inputtomystate_in[14:0], main_inputtomystate_in[24:15], main_inputtomystate_in[24:15], main_inputtomystate_in[14:0]};
  assign zll_main_inputtomystate18_in = {zll_main_inputtomystate_in[49:35], zll_main_inputtomystate_in[34:25], zll_main_inputtomystate_in[34:25], zll_main_inputtomystate_in[49:35]};
  assign zll_main_inputtomystate17_in = {zll_main_inputtomystate18_in[49:35], zll_main_inputtomystate18_in[34:25], zll_main_inputtomystate18_in[34:25], zll_main_inputtomystate18_in[49:35]};
  assign zll_main_inputtomystate9_in = {zll_main_inputtomystate17_in[49:35], zll_main_inputtomystate17_in[34:25], zll_main_inputtomystate17_in[34:25], zll_main_inputtomystate17_in[49:35]};
  assign zll_main_inputtomystate1_in = {zll_main_inputtomystate9_in[34:25], zll_main_inputtomystate9_in[49:35]};
  assign zll_main_inputtomystate3_in = zll_main_inputtomystate1_in[24:0];
  assign zll_main_inputtomystate12_in = {zll_main_inputtomystate3_in[13:9], zll_main_inputtomystate3_in[8:0]};
  assign zll_main_inputtomystate14_in = zll_main_inputtomystate9_in[24:0];
  assign zll_main_inputtomystate13_in = zll_main_inputtomystate17_in[24:0];
  assign zll_main_inputtomystate8_in = {zll_main_inputtomystate13_in[12:9], zll_main_inputtomystate13_in[8:0]};
  assign zll_main_inputtomystate16_in = zll_main_inputtomystate18_in[24:0];
  assign zll_main_inputtomystate2_in = {zll_main_inputtomystate16_in[22:15], zll_main_inputtomystate16_in[14], zll_main_inputtomystate16_in[13:9], zll_main_inputtomystate16_in[8:0]};
  assign zll_main_inputtomystate10_in = zll_main_inputtomystate_in[24:0];
  assign zll_main_inputtomystate11_in = {zll_main_inputtomystate10_in[18:15], zll_main_inputtomystate10_in[14], zll_main_inputtomystate10_in[13:9], zll_main_inputtomystate10_in[8:0]};
  assign zll_main_inputtomystate15_in = {zll_main_inputtomystate11_in[18:15], zll_main_inputtomystate11_in[14], zll_main_inputtomystate11_in[8:0]};
  assign zll_main_incrpipeline5_in = {(zll_main_inputtomystate10_in[24:23] == 2'h0) ? {zll_main_inputtomystate15_in[9], 1'h1, zll_main_inputtomystate15_in[13:10], 5'h0, zll_main_inputtomystate15_in[13:10]} : ((zll_main_inputtomystate16_in[24:23] == 2'h1) ? {zll_main_inputtomystate2_in[14], zll_main_inputtomystate2_in[13:9], 1'h1, zll_main_inputtomystate2_in[22:15]} : (((zll_main_inputtomystate13_in[24:23] == 2'h2) && ((zll_main_inputtomystate13_in[15] == 1'h1) && (zll_main_inputtomystate13_in[13] == 1'h1))) ? {11'h400, zll_main_inputtomystate8_in[12:9]} : (((zll_main_inputtomystate14_in[24:23] == 2'h2) && ((zll_main_inputtomystate14_in[15] == 1'h1) && (zll_main_inputtomystate14_in[13] == 1'h0))) ? {6'h20, zll_main_inputtomystate14_in[8:0]} : {6'h0, zll_main_inputtomystate12_in[8:0]}))), zll_main_loop6_in[29:0]};
  assign zll_main_incrpipeline4_in = zll_main_incrpipeline5_in[44:0];
  assign id_inR1 = zll_main_incrpipeline4_in[29:0];
  assign zll_main_incrpipeline8_in = {zll_main_incrpipeline4_in[44:30], id_inR1[29:15]};
  assign zll_main_incrpipeline6_in = {zll_main_incrpipeline8_in[29:15], zll_main_incrpipeline8_in[14:0]};
  assign id_inR2 = zll_main_incrpipeline6_in[29:0];
  assign zll_main_incrpipeline10_in = zll_main_incrpipeline4_in[29:0];
  assign resize_in = zll_main_incrpipeline10_in[29:0];
  assign binop_in = {128'(resize_in[29:0]), {8'h80{1'h0}}};
  assign resize_inR1 = binop_in[255:128] >> binop_in[127:0];
  assign zll_main_loop1_in = {{id_inR2[29:15], id_inR2[14:0]}, resize_inR1[14:0]};
  assign zll_main_loop4_in = zll_main_loop1_in[44:0];
  assign main_mystatetooutput_in = zll_main_loop4_in[14:0];
  assign zll_main_mystatetooutput4_in = {main_mystatetooutput_in[14:0], main_mystatetooutput_in[14:0]};
  assign zll_main_mystatetooutput7_in = {zll_main_mystatetooutput4_in[29:15], zll_main_mystatetooutput4_in[29:15]};
  assign zll_main_mystatetooutput1_in = zll_main_mystatetooutput7_in[29:15];
  assign zll_main_mystatetooutput3_in = zll_main_mystatetooutput1_in[14:0];
  assign zll_main_mystatetooutput_in = zll_main_mystatetooutput3_in[8:0];
  assign zll_main_mystatetooutput2_in = zll_main_mystatetooutput7_in[14:0];
  assign zll_main_mystatetooutput8_in = {zll_main_mystatetooutput2_in[13:9], zll_main_mystatetooutput2_in[7:0]};
  assign zll_main_mystatetooutput5_in = zll_main_mystatetooutput4_in[14:0];
  assign zll_main_mystatetooutput6_in = {zll_main_mystatetooutput5_in[13:9], zll_main_mystatetooutput5_in[3:0]};
  assign zll_rewire_monad_iterst27_in = {{((zll_main_mystatetooutput5_in[14] == 1'h1) && (zll_main_mystatetooutput5_in[8] == 1'h0)) ? {2'h3, zll_main_mystatetooutput6_in[8:4], 5'h0, zll_main_mystatetooutput6_in[3:0]} : (((zll_main_mystatetooutput2_in[14] == 1'h1) && (zll_main_mystatetooutput2_in[8] == 1'h1)) ? {2'h1, zll_main_mystatetooutput8_in[12:8], 1'h1, zll_main_mystatetooutput8_in[7:0]} : {7'h0, zll_main_mystatetooutput_in[8:0]}), zll_main_loop4_in[44:15]}, zll_rewire_monad_iterst32_in[29:0]};
  assign zll_rewire_monad_iterst25_in = zll_rewire_monad_iterst27_in[75:0];
  assign zll_rewire_monad_iterst36_in = {2'h0, zll_rewire_monad_iterst25_in[75:30], zll_rewire_monad_iterst25_in[29:0]};
  assign zll_rewire_monad_iterst26_in = zll_rewire_monad_iterst36_in[77:0];
  assign zll_rewire_monad_iterst35_in = {zll_rewire_monad_iterst26_in[75:30], zll_rewire_monad_iterst26_in[29:0]};
  assign zll_rewire_monad_iterst22_in = {zll_rewire_monad_iterst35_in[29:0], zll_rewire_monad_iterst35_in[75:30]};
  assign zll_rewire_monad_iterst37_in = {zll_rewire_monad_iterst22_in[45:30], zll_rewire_monad_iterst22_in[75:46], zll_rewire_monad_iterst22_in[29:0]};
  assign zll_rewire_monad_iterst31_in = {zll_rewire_monad_iterst37_in[75:60], zll_rewire_monad_iterst37_in[29:0], zll_rewire_monad_iterst37_in[59:30]};
  assign zll_rewire_monad_iterst15_in = zll_rewire_monad_iterst31_in[59:30];
  assign zll_rewire_monad_iterst4_in = {zll_rewire_monad_iterst31_in[75:60], {{2'h1, {6'h2e{1'h0}}}, zll_rewire_monad_iterst15_in[29:0]}};
  assign zll_rewire_monad_iterst29_in = {zll_rewire_monad_iterst4_in[93:78], zll_rewire_monad_iterst4_in[77:0]};
  assign zll_rewire_monad_iterst33_in = {zll_rewire_monad_iterst29_in[93:78], zll_rewire_monad_iterst29_in[29:0]};
  assign {__padding, __out0, __st0_next} = {{1'h1, {5'h1f{1'h0}}}, zll_rewire_monad_iterst33_in[45:30], zll_rewire_monad_iterst33_in[29:0]};
  initial __st0 = 30'h0;
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      __st0 <= 30'h0;
    end else begin
      __st0 <= __st0_next;
    end
  end
endmodule