module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [99:0] __in0,
  output logic [99:0] __out0,
  output logic [99:0] __out1,
  output logic [99:0] __out2,
  output logic [99:0] __out3);
  logic [99:0] main_dev_in;
  logic [106:0] zll_main_dev2_in;
  logic [0:0] zll_main_dev2_out;
  logic [106:0] zll_main_dev2_inR1;
  logic [0:0] zll_main_dev2_outR1;
  logic [106:0] zll_main_dev2_inR2;
  logic [0:0] zll_main_dev2_outR2;
  logic [106:0] zll_main_dev2_inR3;
  logic [0:0] zll_main_dev2_outR3;
  logic [106:0] zll_main_dev2_inR4;
  logic [0:0] zll_main_dev2_outR4;
  logic [106:0] zll_main_dev2_inR5;
  logic [0:0] zll_main_dev2_outR5;
  logic [106:0] zll_main_dev2_inR6;
  logic [0:0] zll_main_dev2_outR6;
  logic [106:0] zll_main_dev2_inR7;
  logic [0:0] zll_main_dev2_outR7;
  logic [106:0] zll_main_dev2_inR8;
  logic [0:0] zll_main_dev2_outR8;
  logic [106:0] zll_main_dev2_inR9;
  logic [0:0] zll_main_dev2_outR9;
  logic [106:0] zll_main_dev2_inR10;
  logic [0:0] zll_main_dev2_outR10;
  logic [106:0] zll_main_dev2_inR11;
  logic [0:0] zll_main_dev2_outR11;
  logic [106:0] zll_main_dev2_inR12;
  logic [0:0] zll_main_dev2_outR12;
  logic [106:0] zll_main_dev2_inR13;
  logic [0:0] zll_main_dev2_outR13;
  logic [106:0] zll_main_dev2_inR14;
  logic [0:0] zll_main_dev2_outR14;
  logic [106:0] zll_main_dev2_inR15;
  logic [0:0] zll_main_dev2_outR15;
  logic [106:0] zll_main_dev2_inR16;
  logic [0:0] zll_main_dev2_outR16;
  logic [106:0] zll_main_dev2_inR17;
  logic [0:0] zll_main_dev2_outR17;
  logic [106:0] zll_main_dev2_inR18;
  logic [0:0] zll_main_dev2_outR18;
  logic [106:0] zll_main_dev2_inR19;
  logic [0:0] zll_main_dev2_outR19;
  logic [106:0] zll_main_dev2_inR20;
  logic [0:0] zll_main_dev2_outR20;
  logic [106:0] zll_main_dev2_inR21;
  logic [0:0] zll_main_dev2_outR21;
  logic [106:0] zll_main_dev2_inR22;
  logic [0:0] zll_main_dev2_outR22;
  logic [106:0] zll_main_dev2_inR23;
  logic [0:0] zll_main_dev2_outR23;
  logic [106:0] zll_main_dev2_inR24;
  logic [0:0] zll_main_dev2_outR24;
  logic [106:0] zll_main_dev2_inR25;
  logic [0:0] zll_main_dev2_outR25;
  logic [106:0] zll_main_dev2_inR26;
  logic [0:0] zll_main_dev2_outR26;
  logic [106:0] zll_main_dev2_inR27;
  logic [0:0] zll_main_dev2_outR27;
  logic [106:0] zll_main_dev2_inR28;
  logic [0:0] zll_main_dev2_outR28;
  logic [106:0] zll_main_dev2_inR29;
  logic [0:0] zll_main_dev2_outR29;
  logic [106:0] zll_main_dev2_inR30;
  logic [0:0] zll_main_dev2_outR30;
  logic [106:0] zll_main_dev2_inR31;
  logic [0:0] zll_main_dev2_outR31;
  logic [106:0] zll_main_dev2_inR32;
  logic [0:0] zll_main_dev2_outR32;
  logic [106:0] zll_main_dev2_inR33;
  logic [0:0] zll_main_dev2_outR33;
  logic [106:0] zll_main_dev2_inR34;
  logic [0:0] zll_main_dev2_outR34;
  logic [106:0] zll_main_dev2_inR35;
  logic [0:0] zll_main_dev2_outR35;
  logic [106:0] zll_main_dev2_inR36;
  logic [0:0] zll_main_dev2_outR36;
  logic [106:0] zll_main_dev2_inR37;
  logic [0:0] zll_main_dev2_outR37;
  logic [106:0] zll_main_dev2_inR38;
  logic [0:0] zll_main_dev2_outR38;
  logic [106:0] zll_main_dev2_inR39;
  logic [0:0] zll_main_dev2_outR39;
  logic [106:0] zll_main_dev2_inR40;
  logic [0:0] zll_main_dev2_outR40;
  logic [106:0] zll_main_dev2_inR41;
  logic [0:0] zll_main_dev2_outR41;
  logic [106:0] zll_main_dev2_inR42;
  logic [0:0] zll_main_dev2_outR42;
  logic [106:0] zll_main_dev2_inR43;
  logic [0:0] zll_main_dev2_outR43;
  logic [106:0] zll_main_dev2_inR44;
  logic [0:0] zll_main_dev2_outR44;
  logic [106:0] zll_main_dev2_inR45;
  logic [0:0] zll_main_dev2_outR45;
  logic [106:0] zll_main_dev2_inR46;
  logic [0:0] zll_main_dev2_outR46;
  logic [106:0] zll_main_dev2_inR47;
  logic [0:0] zll_main_dev2_outR47;
  logic [106:0] zll_main_dev2_inR48;
  logic [0:0] zll_main_dev2_outR48;
  logic [106:0] zll_main_dev2_inR49;
  logic [0:0] zll_main_dev2_outR49;
  logic [106:0] zll_main_dev2_inR50;
  logic [0:0] zll_main_dev2_outR50;
  logic [106:0] zll_main_dev2_inR51;
  logic [0:0] zll_main_dev2_outR51;
  logic [106:0] zll_main_dev2_inR52;
  logic [0:0] zll_main_dev2_outR52;
  logic [106:0] zll_main_dev2_inR53;
  logic [0:0] zll_main_dev2_outR53;
  logic [106:0] zll_main_dev2_inR54;
  logic [0:0] zll_main_dev2_outR54;
  logic [106:0] zll_main_dev2_inR55;
  logic [0:0] zll_main_dev2_outR55;
  logic [106:0] zll_main_dev2_inR56;
  logic [0:0] zll_main_dev2_outR56;
  logic [106:0] zll_main_dev2_inR57;
  logic [0:0] zll_main_dev2_outR57;
  logic [106:0] zll_main_dev2_inR58;
  logic [0:0] zll_main_dev2_outR58;
  logic [106:0] zll_main_dev2_inR59;
  logic [0:0] zll_main_dev2_outR59;
  logic [106:0] zll_main_dev2_inR60;
  logic [0:0] zll_main_dev2_outR60;
  logic [106:0] zll_main_dev2_inR61;
  logic [0:0] zll_main_dev2_outR61;
  logic [106:0] zll_main_dev2_inR62;
  logic [0:0] zll_main_dev2_outR62;
  logic [106:0] zll_main_dev2_inR63;
  logic [0:0] zll_main_dev2_outR63;
  logic [106:0] zll_main_dev2_inR64;
  logic [0:0] zll_main_dev2_outR64;
  logic [106:0] zll_main_dev2_inR65;
  logic [0:0] zll_main_dev2_outR65;
  logic [106:0] zll_main_dev2_inR66;
  logic [0:0] zll_main_dev2_outR66;
  logic [106:0] zll_main_dev2_inR67;
  logic [0:0] zll_main_dev2_outR67;
  logic [106:0] zll_main_dev2_inR68;
  logic [0:0] zll_main_dev2_outR68;
  logic [106:0] zll_main_dev2_inR69;
  logic [0:0] zll_main_dev2_outR69;
  logic [106:0] zll_main_dev2_inR70;
  logic [0:0] zll_main_dev2_outR70;
  logic [106:0] zll_main_dev2_inR71;
  logic [0:0] zll_main_dev2_outR71;
  logic [106:0] zll_main_dev2_inR72;
  logic [0:0] zll_main_dev2_outR72;
  logic [106:0] zll_main_dev2_inR73;
  logic [0:0] zll_main_dev2_outR73;
  logic [106:0] zll_main_dev2_inR74;
  logic [0:0] zll_main_dev2_outR74;
  logic [106:0] zll_main_dev2_inR75;
  logic [0:0] zll_main_dev2_outR75;
  logic [106:0] zll_main_dev2_inR76;
  logic [0:0] zll_main_dev2_outR76;
  logic [106:0] zll_main_dev2_inR77;
  logic [0:0] zll_main_dev2_outR77;
  logic [106:0] zll_main_dev2_inR78;
  logic [0:0] zll_main_dev2_outR78;
  logic [106:0] zll_main_dev2_inR79;
  logic [0:0] zll_main_dev2_outR79;
  logic [106:0] zll_main_dev2_inR80;
  logic [0:0] zll_main_dev2_outR80;
  logic [106:0] zll_main_dev2_inR81;
  logic [0:0] zll_main_dev2_outR81;
  logic [106:0] zll_main_dev2_inR82;
  logic [0:0] zll_main_dev2_outR82;
  logic [106:0] zll_main_dev2_inR83;
  logic [0:0] zll_main_dev2_outR83;
  logic [106:0] zll_main_dev2_inR84;
  logic [0:0] zll_main_dev2_outR84;
  logic [106:0] zll_main_dev2_inR85;
  logic [0:0] zll_main_dev2_outR85;
  logic [106:0] zll_main_dev2_inR86;
  logic [0:0] zll_main_dev2_outR86;
  logic [106:0] zll_main_dev2_inR87;
  logic [0:0] zll_main_dev2_outR87;
  logic [106:0] zll_main_dev2_inR88;
  logic [0:0] zll_main_dev2_outR88;
  logic [106:0] zll_main_dev2_inR89;
  logic [0:0] zll_main_dev2_outR89;
  logic [106:0] zll_main_dev2_inR90;
  logic [0:0] zll_main_dev2_outR90;
  logic [106:0] zll_main_dev2_inR91;
  logic [0:0] zll_main_dev2_outR91;
  logic [106:0] zll_main_dev2_inR92;
  logic [0:0] zll_main_dev2_outR92;
  logic [106:0] zll_main_dev2_inR93;
  logic [0:0] zll_main_dev2_outR93;
  logic [106:0] zll_main_dev2_inR94;
  logic [0:0] zll_main_dev2_outR94;
  logic [106:0] zll_main_dev2_inR95;
  logic [0:0] zll_main_dev2_outR95;
  logic [106:0] zll_main_dev2_inR96;
  logic [0:0] zll_main_dev2_outR96;
  logic [106:0] zll_main_dev2_inR97;
  logic [0:0] zll_main_dev2_outR97;
  logic [106:0] zll_main_dev2_inR98;
  logic [0:0] zll_main_dev2_outR98;
  logic [106:0] zll_main_dev2_inR99;
  logic [0:0] zll_main_dev2_outR99;
  logic [106:0] zll_main_dev5_in;
  logic [0:0] zll_main_dev5_out;
  logic [106:0] zll_main_dev5_inR1;
  logic [0:0] zll_main_dev5_outR1;
  logic [106:0] zll_main_dev5_inR2;
  logic [0:0] zll_main_dev5_outR2;
  logic [106:0] zll_main_dev5_inR3;
  logic [0:0] zll_main_dev5_outR3;
  logic [106:0] zll_main_dev5_inR4;
  logic [0:0] zll_main_dev5_outR4;
  logic [106:0] zll_main_dev5_inR5;
  logic [0:0] zll_main_dev5_outR5;
  logic [106:0] zll_main_dev5_inR6;
  logic [0:0] zll_main_dev5_outR6;
  logic [106:0] zll_main_dev5_inR7;
  logic [0:0] zll_main_dev5_outR7;
  logic [106:0] zll_main_dev5_inR8;
  logic [0:0] zll_main_dev5_outR8;
  logic [106:0] zll_main_dev5_inR9;
  logic [0:0] zll_main_dev5_outR9;
  logic [106:0] zll_main_dev5_inR10;
  logic [0:0] zll_main_dev5_outR10;
  logic [106:0] zll_main_dev5_inR11;
  logic [0:0] zll_main_dev5_outR11;
  logic [106:0] zll_main_dev5_inR12;
  logic [0:0] zll_main_dev5_outR12;
  logic [106:0] zll_main_dev5_inR13;
  logic [0:0] zll_main_dev5_outR13;
  logic [106:0] zll_main_dev5_inR14;
  logic [0:0] zll_main_dev5_outR14;
  logic [106:0] zll_main_dev5_inR15;
  logic [0:0] zll_main_dev5_outR15;
  logic [106:0] zll_main_dev5_inR16;
  logic [0:0] zll_main_dev5_outR16;
  logic [106:0] zll_main_dev5_inR17;
  logic [0:0] zll_main_dev5_outR17;
  logic [106:0] zll_main_dev5_inR18;
  logic [0:0] zll_main_dev5_outR18;
  logic [106:0] zll_main_dev5_inR19;
  logic [0:0] zll_main_dev5_outR19;
  logic [106:0] zll_main_dev5_inR20;
  logic [0:0] zll_main_dev5_outR20;
  logic [106:0] zll_main_dev5_inR21;
  logic [0:0] zll_main_dev5_outR21;
  logic [106:0] zll_main_dev5_inR22;
  logic [0:0] zll_main_dev5_outR22;
  logic [106:0] zll_main_dev5_inR23;
  logic [0:0] zll_main_dev5_outR23;
  logic [106:0] zll_main_dev5_inR24;
  logic [0:0] zll_main_dev5_outR24;
  logic [106:0] zll_main_dev5_inR25;
  logic [0:0] zll_main_dev5_outR25;
  logic [106:0] zll_main_dev5_inR26;
  logic [0:0] zll_main_dev5_outR26;
  logic [106:0] zll_main_dev5_inR27;
  logic [0:0] zll_main_dev5_outR27;
  logic [106:0] zll_main_dev5_inR28;
  logic [0:0] zll_main_dev5_outR28;
  logic [106:0] zll_main_dev5_inR29;
  logic [0:0] zll_main_dev5_outR29;
  logic [106:0] zll_main_dev5_inR30;
  logic [0:0] zll_main_dev5_outR30;
  logic [106:0] zll_main_dev5_inR31;
  logic [0:0] zll_main_dev5_outR31;
  logic [106:0] zll_main_dev5_inR32;
  logic [0:0] zll_main_dev5_outR32;
  logic [106:0] zll_main_dev5_inR33;
  logic [0:0] zll_main_dev5_outR33;
  logic [106:0] zll_main_dev5_inR34;
  logic [0:0] zll_main_dev5_outR34;
  logic [106:0] zll_main_dev5_inR35;
  logic [0:0] zll_main_dev5_outR35;
  logic [106:0] zll_main_dev5_inR36;
  logic [0:0] zll_main_dev5_outR36;
  logic [106:0] zll_main_dev5_inR37;
  logic [0:0] zll_main_dev5_outR37;
  logic [106:0] zll_main_dev5_inR38;
  logic [0:0] zll_main_dev5_outR38;
  logic [106:0] zll_main_dev5_inR39;
  logic [0:0] zll_main_dev5_outR39;
  logic [106:0] zll_main_dev5_inR40;
  logic [0:0] zll_main_dev5_outR40;
  logic [106:0] zll_main_dev5_inR41;
  logic [0:0] zll_main_dev5_outR41;
  logic [106:0] zll_main_dev5_inR42;
  logic [0:0] zll_main_dev5_outR42;
  logic [106:0] zll_main_dev5_inR43;
  logic [0:0] zll_main_dev5_outR43;
  logic [106:0] zll_main_dev5_inR44;
  logic [0:0] zll_main_dev5_outR44;
  logic [106:0] zll_main_dev5_inR45;
  logic [0:0] zll_main_dev5_outR45;
  logic [106:0] zll_main_dev5_inR46;
  logic [0:0] zll_main_dev5_outR46;
  logic [106:0] zll_main_dev5_inR47;
  logic [0:0] zll_main_dev5_outR47;
  logic [106:0] zll_main_dev5_inR48;
  logic [0:0] zll_main_dev5_outR48;
  logic [106:0] zll_main_dev5_inR49;
  logic [0:0] zll_main_dev5_outR49;
  logic [106:0] zll_main_dev5_inR50;
  logic [0:0] zll_main_dev5_outR50;
  logic [106:0] zll_main_dev5_inR51;
  logic [0:0] zll_main_dev5_outR51;
  logic [106:0] zll_main_dev5_inR52;
  logic [0:0] zll_main_dev5_outR52;
  logic [106:0] zll_main_dev5_inR53;
  logic [0:0] zll_main_dev5_outR53;
  logic [106:0] zll_main_dev5_inR54;
  logic [0:0] zll_main_dev5_outR54;
  logic [106:0] zll_main_dev5_inR55;
  logic [0:0] zll_main_dev5_outR55;
  logic [106:0] zll_main_dev5_inR56;
  logic [0:0] zll_main_dev5_outR56;
  logic [106:0] zll_main_dev5_inR57;
  logic [0:0] zll_main_dev5_outR57;
  logic [106:0] zll_main_dev5_inR58;
  logic [0:0] zll_main_dev5_outR58;
  logic [106:0] zll_main_dev5_inR59;
  logic [0:0] zll_main_dev5_outR59;
  logic [106:0] zll_main_dev5_inR60;
  logic [0:0] zll_main_dev5_outR60;
  logic [106:0] zll_main_dev5_inR61;
  logic [0:0] zll_main_dev5_outR61;
  logic [106:0] zll_main_dev5_inR62;
  logic [0:0] zll_main_dev5_outR62;
  logic [106:0] zll_main_dev5_inR63;
  logic [0:0] zll_main_dev5_outR63;
  logic [106:0] zll_main_dev5_inR64;
  logic [0:0] zll_main_dev5_outR64;
  logic [106:0] zll_main_dev5_inR65;
  logic [0:0] zll_main_dev5_outR65;
  logic [106:0] zll_main_dev5_inR66;
  logic [0:0] zll_main_dev5_outR66;
  logic [106:0] zll_main_dev5_inR67;
  logic [0:0] zll_main_dev5_outR67;
  logic [106:0] zll_main_dev5_inR68;
  logic [0:0] zll_main_dev5_outR68;
  logic [106:0] zll_main_dev5_inR69;
  logic [0:0] zll_main_dev5_outR69;
  logic [106:0] zll_main_dev5_inR70;
  logic [0:0] zll_main_dev5_outR70;
  logic [106:0] zll_main_dev5_inR71;
  logic [0:0] zll_main_dev5_outR71;
  logic [106:0] zll_main_dev5_inR72;
  logic [0:0] zll_main_dev5_outR72;
  logic [106:0] zll_main_dev5_inR73;
  logic [0:0] zll_main_dev5_outR73;
  logic [106:0] zll_main_dev5_inR74;
  logic [0:0] zll_main_dev5_outR74;
  logic [106:0] zll_main_dev5_inR75;
  logic [0:0] zll_main_dev5_outR75;
  logic [106:0] zll_main_dev5_inR76;
  logic [0:0] zll_main_dev5_outR76;
  logic [106:0] zll_main_dev5_inR77;
  logic [0:0] zll_main_dev5_outR77;
  logic [106:0] zll_main_dev5_inR78;
  logic [0:0] zll_main_dev5_outR78;
  logic [106:0] zll_main_dev5_inR79;
  logic [0:0] zll_main_dev5_outR79;
  logic [106:0] zll_main_dev5_inR80;
  logic [0:0] zll_main_dev5_outR80;
  logic [106:0] zll_main_dev5_inR81;
  logic [0:0] zll_main_dev5_outR81;
  logic [106:0] zll_main_dev5_inR82;
  logic [0:0] zll_main_dev5_outR82;
  logic [106:0] zll_main_dev5_inR83;
  logic [0:0] zll_main_dev5_outR83;
  logic [106:0] zll_main_dev5_inR84;
  logic [0:0] zll_main_dev5_outR84;
  logic [106:0] zll_main_dev5_inR85;
  logic [0:0] zll_main_dev5_outR85;
  logic [106:0] zll_main_dev5_inR86;
  logic [0:0] zll_main_dev5_outR86;
  logic [106:0] zll_main_dev5_inR87;
  logic [0:0] zll_main_dev5_outR87;
  logic [106:0] zll_main_dev5_inR88;
  logic [0:0] zll_main_dev5_outR88;
  logic [106:0] zll_main_dev5_inR89;
  logic [0:0] zll_main_dev5_outR89;
  logic [106:0] zll_main_dev5_inR90;
  logic [0:0] zll_main_dev5_outR90;
  logic [106:0] zll_main_dev5_inR91;
  logic [0:0] zll_main_dev5_outR91;
  logic [106:0] zll_main_dev5_inR92;
  logic [0:0] zll_main_dev5_outR92;
  logic [106:0] zll_main_dev5_inR93;
  logic [0:0] zll_main_dev5_outR93;
  logic [106:0] zll_main_dev5_inR94;
  logic [0:0] zll_main_dev5_outR94;
  logic [106:0] zll_main_dev5_inR95;
  logic [0:0] zll_main_dev5_outR95;
  logic [106:0] zll_main_dev5_inR96;
  logic [0:0] zll_main_dev5_outR96;
  logic [106:0] zll_main_dev5_inR97;
  logic [0:0] zll_main_dev5_outR97;
  logic [106:0] zll_main_dev5_inR98;
  logic [0:0] zll_main_dev5_outR98;
  logic [106:0] zll_main_dev5_inR99;
  logic [0:0] zll_main_dev5_outR99;
  logic [106:0] zll_main_dev8_in;
  logic [0:0] zll_main_dev8_out;
  logic [106:0] zll_main_dev8_inR1;
  logic [0:0] zll_main_dev8_outR1;
  logic [106:0] zll_main_dev8_inR2;
  logic [0:0] zll_main_dev8_outR2;
  logic [106:0] zll_main_dev8_inR3;
  logic [0:0] zll_main_dev8_outR3;
  logic [106:0] zll_main_dev8_inR4;
  logic [0:0] zll_main_dev8_outR4;
  logic [106:0] zll_main_dev8_inR5;
  logic [0:0] zll_main_dev8_outR5;
  logic [106:0] zll_main_dev8_inR6;
  logic [0:0] zll_main_dev8_outR6;
  logic [106:0] zll_main_dev8_inR7;
  logic [0:0] zll_main_dev8_outR7;
  logic [106:0] zll_main_dev8_inR8;
  logic [0:0] zll_main_dev8_outR8;
  logic [106:0] zll_main_dev8_inR9;
  logic [0:0] zll_main_dev8_outR9;
  logic [106:0] zll_main_dev8_inR10;
  logic [0:0] zll_main_dev8_outR10;
  logic [106:0] zll_main_dev8_inR11;
  logic [0:0] zll_main_dev8_outR11;
  logic [106:0] zll_main_dev8_inR12;
  logic [0:0] zll_main_dev8_outR12;
  logic [106:0] zll_main_dev8_inR13;
  logic [0:0] zll_main_dev8_outR13;
  logic [106:0] zll_main_dev8_inR14;
  logic [0:0] zll_main_dev8_outR14;
  logic [106:0] zll_main_dev8_inR15;
  logic [0:0] zll_main_dev8_outR15;
  logic [106:0] zll_main_dev8_inR16;
  logic [0:0] zll_main_dev8_outR16;
  logic [106:0] zll_main_dev8_inR17;
  logic [0:0] zll_main_dev8_outR17;
  logic [106:0] zll_main_dev8_inR18;
  logic [0:0] zll_main_dev8_outR18;
  logic [106:0] zll_main_dev8_inR19;
  logic [0:0] zll_main_dev8_outR19;
  logic [106:0] zll_main_dev8_inR20;
  logic [0:0] zll_main_dev8_outR20;
  logic [106:0] zll_main_dev8_inR21;
  logic [0:0] zll_main_dev8_outR21;
  logic [106:0] zll_main_dev8_inR22;
  logic [0:0] zll_main_dev8_outR22;
  logic [106:0] zll_main_dev8_inR23;
  logic [0:0] zll_main_dev8_outR23;
  logic [106:0] zll_main_dev8_inR24;
  logic [0:0] zll_main_dev8_outR24;
  logic [106:0] zll_main_dev8_inR25;
  logic [0:0] zll_main_dev8_outR25;
  logic [106:0] zll_main_dev8_inR26;
  logic [0:0] zll_main_dev8_outR26;
  logic [106:0] zll_main_dev8_inR27;
  logic [0:0] zll_main_dev8_outR27;
  logic [106:0] zll_main_dev8_inR28;
  logic [0:0] zll_main_dev8_outR28;
  logic [106:0] zll_main_dev8_inR29;
  logic [0:0] zll_main_dev8_outR29;
  logic [106:0] zll_main_dev8_inR30;
  logic [0:0] zll_main_dev8_outR30;
  logic [106:0] zll_main_dev8_inR31;
  logic [0:0] zll_main_dev8_outR31;
  logic [106:0] zll_main_dev8_inR32;
  logic [0:0] zll_main_dev8_outR32;
  logic [106:0] zll_main_dev8_inR33;
  logic [0:0] zll_main_dev8_outR33;
  logic [106:0] zll_main_dev8_inR34;
  logic [0:0] zll_main_dev8_outR34;
  logic [106:0] zll_main_dev8_inR35;
  logic [0:0] zll_main_dev8_outR35;
  logic [106:0] zll_main_dev8_inR36;
  logic [0:0] zll_main_dev8_outR36;
  logic [106:0] zll_main_dev8_inR37;
  logic [0:0] zll_main_dev8_outR37;
  logic [106:0] zll_main_dev8_inR38;
  logic [0:0] zll_main_dev8_outR38;
  logic [106:0] zll_main_dev8_inR39;
  logic [0:0] zll_main_dev8_outR39;
  logic [106:0] zll_main_dev8_inR40;
  logic [0:0] zll_main_dev8_outR40;
  logic [106:0] zll_main_dev8_inR41;
  logic [0:0] zll_main_dev8_outR41;
  logic [106:0] zll_main_dev8_inR42;
  logic [0:0] zll_main_dev8_outR42;
  logic [106:0] zll_main_dev8_inR43;
  logic [0:0] zll_main_dev8_outR43;
  logic [106:0] zll_main_dev8_inR44;
  logic [0:0] zll_main_dev8_outR44;
  logic [106:0] zll_main_dev8_inR45;
  logic [0:0] zll_main_dev8_outR45;
  logic [106:0] zll_main_dev8_inR46;
  logic [0:0] zll_main_dev8_outR46;
  logic [106:0] zll_main_dev8_inR47;
  logic [0:0] zll_main_dev8_outR47;
  logic [106:0] zll_main_dev8_inR48;
  logic [0:0] zll_main_dev8_outR48;
  logic [106:0] zll_main_dev8_inR49;
  logic [0:0] zll_main_dev8_outR49;
  logic [106:0] zll_main_dev8_inR50;
  logic [0:0] zll_main_dev8_outR50;
  logic [106:0] zll_main_dev8_inR51;
  logic [0:0] zll_main_dev8_outR51;
  logic [106:0] zll_main_dev8_inR52;
  logic [0:0] zll_main_dev8_outR52;
  logic [106:0] zll_main_dev8_inR53;
  logic [0:0] zll_main_dev8_outR53;
  logic [106:0] zll_main_dev8_inR54;
  logic [0:0] zll_main_dev8_outR54;
  logic [106:0] zll_main_dev8_inR55;
  logic [0:0] zll_main_dev8_outR55;
  logic [106:0] zll_main_dev8_inR56;
  logic [0:0] zll_main_dev8_outR56;
  logic [106:0] zll_main_dev8_inR57;
  logic [0:0] zll_main_dev8_outR57;
  logic [106:0] zll_main_dev8_inR58;
  logic [0:0] zll_main_dev8_outR58;
  logic [106:0] zll_main_dev8_inR59;
  logic [0:0] zll_main_dev8_outR59;
  logic [106:0] zll_main_dev8_inR60;
  logic [0:0] zll_main_dev8_outR60;
  logic [106:0] zll_main_dev8_inR61;
  logic [0:0] zll_main_dev8_outR61;
  logic [106:0] zll_main_dev8_inR62;
  logic [0:0] zll_main_dev8_outR62;
  logic [106:0] zll_main_dev8_inR63;
  logic [0:0] zll_main_dev8_outR63;
  logic [106:0] zll_main_dev8_inR64;
  logic [0:0] zll_main_dev8_outR64;
  logic [106:0] zll_main_dev8_inR65;
  logic [0:0] zll_main_dev8_outR65;
  logic [106:0] zll_main_dev8_inR66;
  logic [0:0] zll_main_dev8_outR66;
  logic [106:0] zll_main_dev8_inR67;
  logic [0:0] zll_main_dev8_outR67;
  logic [106:0] zll_main_dev8_inR68;
  logic [0:0] zll_main_dev8_outR68;
  logic [106:0] zll_main_dev8_inR69;
  logic [0:0] zll_main_dev8_outR69;
  logic [106:0] zll_main_dev8_inR70;
  logic [0:0] zll_main_dev8_outR70;
  logic [106:0] zll_main_dev8_inR71;
  logic [0:0] zll_main_dev8_outR71;
  logic [106:0] zll_main_dev8_inR72;
  logic [0:0] zll_main_dev8_outR72;
  logic [106:0] zll_main_dev8_inR73;
  logic [0:0] zll_main_dev8_outR73;
  logic [106:0] zll_main_dev8_inR74;
  logic [0:0] zll_main_dev8_outR74;
  logic [106:0] zll_main_dev8_inR75;
  logic [0:0] zll_main_dev8_outR75;
  logic [106:0] zll_main_dev8_inR76;
  logic [0:0] zll_main_dev8_outR76;
  logic [106:0] zll_main_dev8_inR77;
  logic [0:0] zll_main_dev8_outR77;
  logic [106:0] zll_main_dev8_inR78;
  logic [0:0] zll_main_dev8_outR78;
  logic [106:0] zll_main_dev8_inR79;
  logic [0:0] zll_main_dev8_outR79;
  logic [106:0] zll_main_dev8_inR80;
  logic [0:0] zll_main_dev8_outR80;
  logic [106:0] zll_main_dev8_inR81;
  logic [0:0] zll_main_dev8_outR81;
  logic [106:0] zll_main_dev8_inR82;
  logic [0:0] zll_main_dev8_outR82;
  logic [106:0] zll_main_dev8_inR83;
  logic [0:0] zll_main_dev8_outR83;
  logic [106:0] zll_main_dev8_inR84;
  logic [0:0] zll_main_dev8_outR84;
  logic [106:0] zll_main_dev8_inR85;
  logic [0:0] zll_main_dev8_outR85;
  logic [106:0] zll_main_dev8_inR86;
  logic [0:0] zll_main_dev8_outR86;
  logic [106:0] zll_main_dev8_inR87;
  logic [0:0] zll_main_dev8_outR87;
  logic [106:0] zll_main_dev8_inR88;
  logic [0:0] zll_main_dev8_outR88;
  logic [106:0] zll_main_dev8_inR89;
  logic [0:0] zll_main_dev8_outR89;
  logic [106:0] zll_main_dev8_inR90;
  logic [0:0] zll_main_dev8_outR90;
  logic [106:0] zll_main_dev8_inR91;
  logic [0:0] zll_main_dev8_outR91;
  logic [106:0] zll_main_dev8_inR92;
  logic [0:0] zll_main_dev8_outR92;
  logic [106:0] zll_main_dev8_inR93;
  logic [0:0] zll_main_dev8_outR93;
  logic [106:0] zll_main_dev8_inR94;
  logic [0:0] zll_main_dev8_outR94;
  logic [106:0] zll_main_dev8_inR95;
  logic [0:0] zll_main_dev8_outR95;
  logic [106:0] zll_main_dev8_inR96;
  logic [0:0] zll_main_dev8_outR96;
  logic [106:0] zll_main_dev8_inR97;
  logic [0:0] zll_main_dev8_outR97;
  logic [106:0] zll_main_dev8_inR98;
  logic [0:0] zll_main_dev8_outR98;
  logic [106:0] zll_main_dev8_inR99;
  logic [0:0] zll_main_dev8_outR99;
  logic [106:0] zll_main_dev11_in;
  logic [0:0] zll_main_dev11_out;
  logic [106:0] zll_main_dev11_inR1;
  logic [0:0] zll_main_dev11_outR1;
  logic [106:0] zll_main_dev11_inR2;
  logic [0:0] zll_main_dev11_outR2;
  logic [106:0] zll_main_dev11_inR3;
  logic [0:0] zll_main_dev11_outR3;
  logic [106:0] zll_main_dev11_inR4;
  logic [0:0] zll_main_dev11_outR4;
  logic [106:0] zll_main_dev11_inR5;
  logic [0:0] zll_main_dev11_outR5;
  logic [106:0] zll_main_dev11_inR6;
  logic [0:0] zll_main_dev11_outR6;
  logic [106:0] zll_main_dev11_inR7;
  logic [0:0] zll_main_dev11_outR7;
  logic [106:0] zll_main_dev11_inR8;
  logic [0:0] zll_main_dev11_outR8;
  logic [106:0] zll_main_dev11_inR9;
  logic [0:0] zll_main_dev11_outR9;
  logic [106:0] zll_main_dev11_inR10;
  logic [0:0] zll_main_dev11_outR10;
  logic [106:0] zll_main_dev11_inR11;
  logic [0:0] zll_main_dev11_outR11;
  logic [106:0] zll_main_dev11_inR12;
  logic [0:0] zll_main_dev11_outR12;
  logic [106:0] zll_main_dev11_inR13;
  logic [0:0] zll_main_dev11_outR13;
  logic [106:0] zll_main_dev11_inR14;
  logic [0:0] zll_main_dev11_outR14;
  logic [106:0] zll_main_dev11_inR15;
  logic [0:0] zll_main_dev11_outR15;
  logic [106:0] zll_main_dev11_inR16;
  logic [0:0] zll_main_dev11_outR16;
  logic [106:0] zll_main_dev11_inR17;
  logic [0:0] zll_main_dev11_outR17;
  logic [106:0] zll_main_dev11_inR18;
  logic [0:0] zll_main_dev11_outR18;
  logic [106:0] zll_main_dev11_inR19;
  logic [0:0] zll_main_dev11_outR19;
  logic [106:0] zll_main_dev11_inR20;
  logic [0:0] zll_main_dev11_outR20;
  logic [106:0] zll_main_dev11_inR21;
  logic [0:0] zll_main_dev11_outR21;
  logic [106:0] zll_main_dev11_inR22;
  logic [0:0] zll_main_dev11_outR22;
  logic [106:0] zll_main_dev11_inR23;
  logic [0:0] zll_main_dev11_outR23;
  logic [106:0] zll_main_dev11_inR24;
  logic [0:0] zll_main_dev11_outR24;
  logic [106:0] zll_main_dev11_inR25;
  logic [0:0] zll_main_dev11_outR25;
  logic [106:0] zll_main_dev11_inR26;
  logic [0:0] zll_main_dev11_outR26;
  logic [106:0] zll_main_dev11_inR27;
  logic [0:0] zll_main_dev11_outR27;
  logic [106:0] zll_main_dev11_inR28;
  logic [0:0] zll_main_dev11_outR28;
  logic [106:0] zll_main_dev11_inR29;
  logic [0:0] zll_main_dev11_outR29;
  logic [106:0] zll_main_dev11_inR30;
  logic [0:0] zll_main_dev11_outR30;
  logic [106:0] zll_main_dev11_inR31;
  logic [0:0] zll_main_dev11_outR31;
  logic [106:0] zll_main_dev11_inR32;
  logic [0:0] zll_main_dev11_outR32;
  logic [106:0] zll_main_dev11_inR33;
  logic [0:0] zll_main_dev11_outR33;
  logic [106:0] zll_main_dev11_inR34;
  logic [0:0] zll_main_dev11_outR34;
  logic [106:0] zll_main_dev11_inR35;
  logic [0:0] zll_main_dev11_outR35;
  logic [106:0] zll_main_dev11_inR36;
  logic [0:0] zll_main_dev11_outR36;
  logic [106:0] zll_main_dev11_inR37;
  logic [0:0] zll_main_dev11_outR37;
  logic [106:0] zll_main_dev11_inR38;
  logic [0:0] zll_main_dev11_outR38;
  logic [106:0] zll_main_dev11_inR39;
  logic [0:0] zll_main_dev11_outR39;
  logic [106:0] zll_main_dev11_inR40;
  logic [0:0] zll_main_dev11_outR40;
  logic [106:0] zll_main_dev11_inR41;
  logic [0:0] zll_main_dev11_outR41;
  logic [106:0] zll_main_dev11_inR42;
  logic [0:0] zll_main_dev11_outR42;
  logic [106:0] zll_main_dev11_inR43;
  logic [0:0] zll_main_dev11_outR43;
  logic [106:0] zll_main_dev11_inR44;
  logic [0:0] zll_main_dev11_outR44;
  logic [106:0] zll_main_dev11_inR45;
  logic [0:0] zll_main_dev11_outR45;
  logic [106:0] zll_main_dev11_inR46;
  logic [0:0] zll_main_dev11_outR46;
  logic [106:0] zll_main_dev11_inR47;
  logic [0:0] zll_main_dev11_outR47;
  logic [106:0] zll_main_dev11_inR48;
  logic [0:0] zll_main_dev11_outR48;
  logic [106:0] zll_main_dev11_inR49;
  logic [0:0] zll_main_dev11_outR49;
  logic [106:0] zll_main_dev11_inR50;
  logic [0:0] zll_main_dev11_outR50;
  logic [106:0] zll_main_dev11_inR51;
  logic [0:0] zll_main_dev11_outR51;
  logic [106:0] zll_main_dev11_inR52;
  logic [0:0] zll_main_dev11_outR52;
  logic [106:0] zll_main_dev11_inR53;
  logic [0:0] zll_main_dev11_outR53;
  logic [106:0] zll_main_dev11_inR54;
  logic [0:0] zll_main_dev11_outR54;
  logic [106:0] zll_main_dev11_inR55;
  logic [0:0] zll_main_dev11_outR55;
  logic [106:0] zll_main_dev11_inR56;
  logic [0:0] zll_main_dev11_outR56;
  logic [106:0] zll_main_dev11_inR57;
  logic [0:0] zll_main_dev11_outR57;
  logic [106:0] zll_main_dev11_inR58;
  logic [0:0] zll_main_dev11_outR58;
  logic [106:0] zll_main_dev11_inR59;
  logic [0:0] zll_main_dev11_outR59;
  logic [106:0] zll_main_dev11_inR60;
  logic [0:0] zll_main_dev11_outR60;
  logic [106:0] zll_main_dev11_inR61;
  logic [0:0] zll_main_dev11_outR61;
  logic [106:0] zll_main_dev11_inR62;
  logic [0:0] zll_main_dev11_outR62;
  logic [106:0] zll_main_dev11_inR63;
  logic [0:0] zll_main_dev11_outR63;
  logic [106:0] zll_main_dev11_inR64;
  logic [0:0] zll_main_dev11_outR64;
  logic [106:0] zll_main_dev11_inR65;
  logic [0:0] zll_main_dev11_outR65;
  logic [106:0] zll_main_dev11_inR66;
  logic [0:0] zll_main_dev11_outR66;
  logic [106:0] zll_main_dev11_inR67;
  logic [0:0] zll_main_dev11_outR67;
  logic [106:0] zll_main_dev11_inR68;
  logic [0:0] zll_main_dev11_outR68;
  logic [106:0] zll_main_dev11_inR69;
  logic [0:0] zll_main_dev11_outR69;
  logic [106:0] zll_main_dev11_inR70;
  logic [0:0] zll_main_dev11_outR70;
  logic [106:0] zll_main_dev11_inR71;
  logic [0:0] zll_main_dev11_outR71;
  logic [106:0] zll_main_dev11_inR72;
  logic [0:0] zll_main_dev11_outR72;
  logic [106:0] zll_main_dev11_inR73;
  logic [0:0] zll_main_dev11_outR73;
  logic [106:0] zll_main_dev11_inR74;
  logic [0:0] zll_main_dev11_outR74;
  logic [106:0] zll_main_dev11_inR75;
  logic [0:0] zll_main_dev11_outR75;
  logic [106:0] zll_main_dev11_inR76;
  logic [0:0] zll_main_dev11_outR76;
  logic [106:0] zll_main_dev11_inR77;
  logic [0:0] zll_main_dev11_outR77;
  logic [106:0] zll_main_dev11_inR78;
  logic [0:0] zll_main_dev11_outR78;
  logic [106:0] zll_main_dev11_inR79;
  logic [0:0] zll_main_dev11_outR79;
  logic [106:0] zll_main_dev11_inR80;
  logic [0:0] zll_main_dev11_outR80;
  logic [106:0] zll_main_dev11_inR81;
  logic [0:0] zll_main_dev11_outR81;
  logic [106:0] zll_main_dev11_inR82;
  logic [0:0] zll_main_dev11_outR82;
  logic [106:0] zll_main_dev11_inR83;
  logic [0:0] zll_main_dev11_outR83;
  logic [106:0] zll_main_dev11_inR84;
  logic [0:0] zll_main_dev11_outR84;
  logic [106:0] zll_main_dev11_inR85;
  logic [0:0] zll_main_dev11_outR85;
  logic [106:0] zll_main_dev11_inR86;
  logic [0:0] zll_main_dev11_outR86;
  logic [106:0] zll_main_dev11_inR87;
  logic [0:0] zll_main_dev11_outR87;
  logic [106:0] zll_main_dev11_inR88;
  logic [0:0] zll_main_dev11_outR88;
  logic [106:0] zll_main_dev11_inR89;
  logic [0:0] zll_main_dev11_outR89;
  logic [106:0] zll_main_dev11_inR90;
  logic [0:0] zll_main_dev11_outR90;
  logic [106:0] zll_main_dev11_inR91;
  logic [0:0] zll_main_dev11_outR91;
  logic [106:0] zll_main_dev11_inR92;
  logic [0:0] zll_main_dev11_outR92;
  logic [106:0] zll_main_dev11_inR93;
  logic [0:0] zll_main_dev11_outR93;
  logic [106:0] zll_main_dev11_inR94;
  logic [0:0] zll_main_dev11_outR94;
  logic [106:0] zll_main_dev11_inR95;
  logic [0:0] zll_main_dev11_outR95;
  logic [106:0] zll_main_dev11_inR96;
  logic [0:0] zll_main_dev11_outR96;
  logic [106:0] zll_main_dev11_inR97;
  logic [0:0] zll_main_dev11_outR97;
  logic [106:0] zll_main_dev11_inR98;
  logic [0:0] zll_main_dev11_outR98;
  logic [106:0] zll_main_dev11_inR99;
  logic [0:0] zll_main_dev11_outR99;
  logic [0:0] __continue;
  logic [99:0] __resumption_tag;
  logic [99:0] __resumption_tag_next;
  assign main_dev_in = __resumption_tag;
  assign zll_main_dev2_in = {main_dev_in[99:0], 7'h00};
  ZLL_Main_dev2  inst (zll_main_dev2_in[106:7], zll_main_dev2_in[6:0], zll_main_dev2_out);
  assign zll_main_dev2_inR1 = {main_dev_in[99:0], 7'h01};
  ZLL_Main_dev2  instR1 (zll_main_dev2_inR1[106:7], zll_main_dev2_inR1[6:0], zll_main_dev2_outR1);
  assign zll_main_dev2_inR2 = {main_dev_in[99:0], 7'h02};
  ZLL_Main_dev2  instR2 (zll_main_dev2_inR2[106:7], zll_main_dev2_inR2[6:0], zll_main_dev2_outR2);
  assign zll_main_dev2_inR3 = {main_dev_in[99:0], 7'h03};
  ZLL_Main_dev2  instR3 (zll_main_dev2_inR3[106:7], zll_main_dev2_inR3[6:0], zll_main_dev2_outR3);
  assign zll_main_dev2_inR4 = {main_dev_in[99:0], 7'h04};
  ZLL_Main_dev2  instR4 (zll_main_dev2_inR4[106:7], zll_main_dev2_inR4[6:0], zll_main_dev2_outR4);
  assign zll_main_dev2_inR5 = {main_dev_in[99:0], 7'h05};
  ZLL_Main_dev2  instR5 (zll_main_dev2_inR5[106:7], zll_main_dev2_inR5[6:0], zll_main_dev2_outR5);
  assign zll_main_dev2_inR6 = {main_dev_in[99:0], 7'h06};
  ZLL_Main_dev2  instR6 (zll_main_dev2_inR6[106:7], zll_main_dev2_inR6[6:0], zll_main_dev2_outR6);
  assign zll_main_dev2_inR7 = {main_dev_in[99:0], 7'h07};
  ZLL_Main_dev2  instR7 (zll_main_dev2_inR7[106:7], zll_main_dev2_inR7[6:0], zll_main_dev2_outR7);
  assign zll_main_dev2_inR8 = {main_dev_in[99:0], 7'h08};
  ZLL_Main_dev2  instR8 (zll_main_dev2_inR8[106:7], zll_main_dev2_inR8[6:0], zll_main_dev2_outR8);
  assign zll_main_dev2_inR9 = {main_dev_in[99:0], 7'h09};
  ZLL_Main_dev2  instR9 (zll_main_dev2_inR9[106:7], zll_main_dev2_inR9[6:0], zll_main_dev2_outR9);
  assign zll_main_dev2_inR10 = {main_dev_in[99:0], 7'h0a};
  ZLL_Main_dev2  instR10 (zll_main_dev2_inR10[106:7], zll_main_dev2_inR10[6:0], zll_main_dev2_outR10);
  assign zll_main_dev2_inR11 = {main_dev_in[99:0], 7'h0b};
  ZLL_Main_dev2  instR11 (zll_main_dev2_inR11[106:7], zll_main_dev2_inR11[6:0], zll_main_dev2_outR11);
  assign zll_main_dev2_inR12 = {main_dev_in[99:0], 7'h0c};
  ZLL_Main_dev2  instR12 (zll_main_dev2_inR12[106:7], zll_main_dev2_inR12[6:0], zll_main_dev2_outR12);
  assign zll_main_dev2_inR13 = {main_dev_in[99:0], 7'h0d};
  ZLL_Main_dev2  instR13 (zll_main_dev2_inR13[106:7], zll_main_dev2_inR13[6:0], zll_main_dev2_outR13);
  assign zll_main_dev2_inR14 = {main_dev_in[99:0], 7'h0e};
  ZLL_Main_dev2  instR14 (zll_main_dev2_inR14[106:7], zll_main_dev2_inR14[6:0], zll_main_dev2_outR14);
  assign zll_main_dev2_inR15 = {main_dev_in[99:0], 7'h0f};
  ZLL_Main_dev2  instR15 (zll_main_dev2_inR15[106:7], zll_main_dev2_inR15[6:0], zll_main_dev2_outR15);
  assign zll_main_dev2_inR16 = {main_dev_in[99:0], 7'h10};
  ZLL_Main_dev2  instR16 (zll_main_dev2_inR16[106:7], zll_main_dev2_inR16[6:0], zll_main_dev2_outR16);
  assign zll_main_dev2_inR17 = {main_dev_in[99:0], 7'h11};
  ZLL_Main_dev2  instR17 (zll_main_dev2_inR17[106:7], zll_main_dev2_inR17[6:0], zll_main_dev2_outR17);
  assign zll_main_dev2_inR18 = {main_dev_in[99:0], 7'h12};
  ZLL_Main_dev2  instR18 (zll_main_dev2_inR18[106:7], zll_main_dev2_inR18[6:0], zll_main_dev2_outR18);
  assign zll_main_dev2_inR19 = {main_dev_in[99:0], 7'h13};
  ZLL_Main_dev2  instR19 (zll_main_dev2_inR19[106:7], zll_main_dev2_inR19[6:0], zll_main_dev2_outR19);
  assign zll_main_dev2_inR20 = {main_dev_in[99:0], 7'h14};
  ZLL_Main_dev2  instR20 (zll_main_dev2_inR20[106:7], zll_main_dev2_inR20[6:0], zll_main_dev2_outR20);
  assign zll_main_dev2_inR21 = {main_dev_in[99:0], 7'h15};
  ZLL_Main_dev2  instR21 (zll_main_dev2_inR21[106:7], zll_main_dev2_inR21[6:0], zll_main_dev2_outR21);
  assign zll_main_dev2_inR22 = {main_dev_in[99:0], 7'h16};
  ZLL_Main_dev2  instR22 (zll_main_dev2_inR22[106:7], zll_main_dev2_inR22[6:0], zll_main_dev2_outR22);
  assign zll_main_dev2_inR23 = {main_dev_in[99:0], 7'h17};
  ZLL_Main_dev2  instR23 (zll_main_dev2_inR23[106:7], zll_main_dev2_inR23[6:0], zll_main_dev2_outR23);
  assign zll_main_dev2_inR24 = {main_dev_in[99:0], 7'h18};
  ZLL_Main_dev2  instR24 (zll_main_dev2_inR24[106:7], zll_main_dev2_inR24[6:0], zll_main_dev2_outR24);
  assign zll_main_dev2_inR25 = {main_dev_in[99:0], 7'h19};
  ZLL_Main_dev2  instR25 (zll_main_dev2_inR25[106:7], zll_main_dev2_inR25[6:0], zll_main_dev2_outR25);
  assign zll_main_dev2_inR26 = {main_dev_in[99:0], 7'h1a};
  ZLL_Main_dev2  instR26 (zll_main_dev2_inR26[106:7], zll_main_dev2_inR26[6:0], zll_main_dev2_outR26);
  assign zll_main_dev2_inR27 = {main_dev_in[99:0], 7'h1b};
  ZLL_Main_dev2  instR27 (zll_main_dev2_inR27[106:7], zll_main_dev2_inR27[6:0], zll_main_dev2_outR27);
  assign zll_main_dev2_inR28 = {main_dev_in[99:0], 7'h1c};
  ZLL_Main_dev2  instR28 (zll_main_dev2_inR28[106:7], zll_main_dev2_inR28[6:0], zll_main_dev2_outR28);
  assign zll_main_dev2_inR29 = {main_dev_in[99:0], 7'h1d};
  ZLL_Main_dev2  instR29 (zll_main_dev2_inR29[106:7], zll_main_dev2_inR29[6:0], zll_main_dev2_outR29);
  assign zll_main_dev2_inR30 = {main_dev_in[99:0], 7'h1e};
  ZLL_Main_dev2  instR30 (zll_main_dev2_inR30[106:7], zll_main_dev2_inR30[6:0], zll_main_dev2_outR30);
  assign zll_main_dev2_inR31 = {main_dev_in[99:0], 7'h1f};
  ZLL_Main_dev2  instR31 (zll_main_dev2_inR31[106:7], zll_main_dev2_inR31[6:0], zll_main_dev2_outR31);
  assign zll_main_dev2_inR32 = {main_dev_in[99:0], 7'h20};
  ZLL_Main_dev2  instR32 (zll_main_dev2_inR32[106:7], zll_main_dev2_inR32[6:0], zll_main_dev2_outR32);
  assign zll_main_dev2_inR33 = {main_dev_in[99:0], 7'h21};
  ZLL_Main_dev2  instR33 (zll_main_dev2_inR33[106:7], zll_main_dev2_inR33[6:0], zll_main_dev2_outR33);
  assign zll_main_dev2_inR34 = {main_dev_in[99:0], 7'h22};
  ZLL_Main_dev2  instR34 (zll_main_dev2_inR34[106:7], zll_main_dev2_inR34[6:0], zll_main_dev2_outR34);
  assign zll_main_dev2_inR35 = {main_dev_in[99:0], 7'h23};
  ZLL_Main_dev2  instR35 (zll_main_dev2_inR35[106:7], zll_main_dev2_inR35[6:0], zll_main_dev2_outR35);
  assign zll_main_dev2_inR36 = {main_dev_in[99:0], 7'h24};
  ZLL_Main_dev2  instR36 (zll_main_dev2_inR36[106:7], zll_main_dev2_inR36[6:0], zll_main_dev2_outR36);
  assign zll_main_dev2_inR37 = {main_dev_in[99:0], 7'h25};
  ZLL_Main_dev2  instR37 (zll_main_dev2_inR37[106:7], zll_main_dev2_inR37[6:0], zll_main_dev2_outR37);
  assign zll_main_dev2_inR38 = {main_dev_in[99:0], 7'h26};
  ZLL_Main_dev2  instR38 (zll_main_dev2_inR38[106:7], zll_main_dev2_inR38[6:0], zll_main_dev2_outR38);
  assign zll_main_dev2_inR39 = {main_dev_in[99:0], 7'h27};
  ZLL_Main_dev2  instR39 (zll_main_dev2_inR39[106:7], zll_main_dev2_inR39[6:0], zll_main_dev2_outR39);
  assign zll_main_dev2_inR40 = {main_dev_in[99:0], 7'h28};
  ZLL_Main_dev2  instR40 (zll_main_dev2_inR40[106:7], zll_main_dev2_inR40[6:0], zll_main_dev2_outR40);
  assign zll_main_dev2_inR41 = {main_dev_in[99:0], 7'h29};
  ZLL_Main_dev2  instR41 (zll_main_dev2_inR41[106:7], zll_main_dev2_inR41[6:0], zll_main_dev2_outR41);
  assign zll_main_dev2_inR42 = {main_dev_in[99:0], 7'h2a};
  ZLL_Main_dev2  instR42 (zll_main_dev2_inR42[106:7], zll_main_dev2_inR42[6:0], zll_main_dev2_outR42);
  assign zll_main_dev2_inR43 = {main_dev_in[99:0], 7'h2b};
  ZLL_Main_dev2  instR43 (zll_main_dev2_inR43[106:7], zll_main_dev2_inR43[6:0], zll_main_dev2_outR43);
  assign zll_main_dev2_inR44 = {main_dev_in[99:0], 7'h2c};
  ZLL_Main_dev2  instR44 (zll_main_dev2_inR44[106:7], zll_main_dev2_inR44[6:0], zll_main_dev2_outR44);
  assign zll_main_dev2_inR45 = {main_dev_in[99:0], 7'h2d};
  ZLL_Main_dev2  instR45 (zll_main_dev2_inR45[106:7], zll_main_dev2_inR45[6:0], zll_main_dev2_outR45);
  assign zll_main_dev2_inR46 = {main_dev_in[99:0], 7'h2e};
  ZLL_Main_dev2  instR46 (zll_main_dev2_inR46[106:7], zll_main_dev2_inR46[6:0], zll_main_dev2_outR46);
  assign zll_main_dev2_inR47 = {main_dev_in[99:0], 7'h2f};
  ZLL_Main_dev2  instR47 (zll_main_dev2_inR47[106:7], zll_main_dev2_inR47[6:0], zll_main_dev2_outR47);
  assign zll_main_dev2_inR48 = {main_dev_in[99:0], 7'h30};
  ZLL_Main_dev2  instR48 (zll_main_dev2_inR48[106:7], zll_main_dev2_inR48[6:0], zll_main_dev2_outR48);
  assign zll_main_dev2_inR49 = {main_dev_in[99:0], 7'h31};
  ZLL_Main_dev2  instR49 (zll_main_dev2_inR49[106:7], zll_main_dev2_inR49[6:0], zll_main_dev2_outR49);
  assign zll_main_dev2_inR50 = {main_dev_in[99:0], 7'h32};
  ZLL_Main_dev2  instR50 (zll_main_dev2_inR50[106:7], zll_main_dev2_inR50[6:0], zll_main_dev2_outR50);
  assign zll_main_dev2_inR51 = {main_dev_in[99:0], 7'h33};
  ZLL_Main_dev2  instR51 (zll_main_dev2_inR51[106:7], zll_main_dev2_inR51[6:0], zll_main_dev2_outR51);
  assign zll_main_dev2_inR52 = {main_dev_in[99:0], 7'h34};
  ZLL_Main_dev2  instR52 (zll_main_dev2_inR52[106:7], zll_main_dev2_inR52[6:0], zll_main_dev2_outR52);
  assign zll_main_dev2_inR53 = {main_dev_in[99:0], 7'h35};
  ZLL_Main_dev2  instR53 (zll_main_dev2_inR53[106:7], zll_main_dev2_inR53[6:0], zll_main_dev2_outR53);
  assign zll_main_dev2_inR54 = {main_dev_in[99:0], 7'h36};
  ZLL_Main_dev2  instR54 (zll_main_dev2_inR54[106:7], zll_main_dev2_inR54[6:0], zll_main_dev2_outR54);
  assign zll_main_dev2_inR55 = {main_dev_in[99:0], 7'h37};
  ZLL_Main_dev2  instR55 (zll_main_dev2_inR55[106:7], zll_main_dev2_inR55[6:0], zll_main_dev2_outR55);
  assign zll_main_dev2_inR56 = {main_dev_in[99:0], 7'h38};
  ZLL_Main_dev2  instR56 (zll_main_dev2_inR56[106:7], zll_main_dev2_inR56[6:0], zll_main_dev2_outR56);
  assign zll_main_dev2_inR57 = {main_dev_in[99:0], 7'h39};
  ZLL_Main_dev2  instR57 (zll_main_dev2_inR57[106:7], zll_main_dev2_inR57[6:0], zll_main_dev2_outR57);
  assign zll_main_dev2_inR58 = {main_dev_in[99:0], 7'h3a};
  ZLL_Main_dev2  instR58 (zll_main_dev2_inR58[106:7], zll_main_dev2_inR58[6:0], zll_main_dev2_outR58);
  assign zll_main_dev2_inR59 = {main_dev_in[99:0], 7'h3b};
  ZLL_Main_dev2  instR59 (zll_main_dev2_inR59[106:7], zll_main_dev2_inR59[6:0], zll_main_dev2_outR59);
  assign zll_main_dev2_inR60 = {main_dev_in[99:0], 7'h3c};
  ZLL_Main_dev2  instR60 (zll_main_dev2_inR60[106:7], zll_main_dev2_inR60[6:0], zll_main_dev2_outR60);
  assign zll_main_dev2_inR61 = {main_dev_in[99:0], 7'h3d};
  ZLL_Main_dev2  instR61 (zll_main_dev2_inR61[106:7], zll_main_dev2_inR61[6:0], zll_main_dev2_outR61);
  assign zll_main_dev2_inR62 = {main_dev_in[99:0], 7'h3e};
  ZLL_Main_dev2  instR62 (zll_main_dev2_inR62[106:7], zll_main_dev2_inR62[6:0], zll_main_dev2_outR62);
  assign zll_main_dev2_inR63 = {main_dev_in[99:0], 7'h3f};
  ZLL_Main_dev2  instR63 (zll_main_dev2_inR63[106:7], zll_main_dev2_inR63[6:0], zll_main_dev2_outR63);
  assign zll_main_dev2_inR64 = {main_dev_in[99:0], 7'h40};
  ZLL_Main_dev2  instR64 (zll_main_dev2_inR64[106:7], zll_main_dev2_inR64[6:0], zll_main_dev2_outR64);
  assign zll_main_dev2_inR65 = {main_dev_in[99:0], 7'h41};
  ZLL_Main_dev2  instR65 (zll_main_dev2_inR65[106:7], zll_main_dev2_inR65[6:0], zll_main_dev2_outR65);
  assign zll_main_dev2_inR66 = {main_dev_in[99:0], 7'h42};
  ZLL_Main_dev2  instR66 (zll_main_dev2_inR66[106:7], zll_main_dev2_inR66[6:0], zll_main_dev2_outR66);
  assign zll_main_dev2_inR67 = {main_dev_in[99:0], 7'h43};
  ZLL_Main_dev2  instR67 (zll_main_dev2_inR67[106:7], zll_main_dev2_inR67[6:0], zll_main_dev2_outR67);
  assign zll_main_dev2_inR68 = {main_dev_in[99:0], 7'h44};
  ZLL_Main_dev2  instR68 (zll_main_dev2_inR68[106:7], zll_main_dev2_inR68[6:0], zll_main_dev2_outR68);
  assign zll_main_dev2_inR69 = {main_dev_in[99:0], 7'h45};
  ZLL_Main_dev2  instR69 (zll_main_dev2_inR69[106:7], zll_main_dev2_inR69[6:0], zll_main_dev2_outR69);
  assign zll_main_dev2_inR70 = {main_dev_in[99:0], 7'h46};
  ZLL_Main_dev2  instR70 (zll_main_dev2_inR70[106:7], zll_main_dev2_inR70[6:0], zll_main_dev2_outR70);
  assign zll_main_dev2_inR71 = {main_dev_in[99:0], 7'h47};
  ZLL_Main_dev2  instR71 (zll_main_dev2_inR71[106:7], zll_main_dev2_inR71[6:0], zll_main_dev2_outR71);
  assign zll_main_dev2_inR72 = {main_dev_in[99:0], 7'h48};
  ZLL_Main_dev2  instR72 (zll_main_dev2_inR72[106:7], zll_main_dev2_inR72[6:0], zll_main_dev2_outR72);
  assign zll_main_dev2_inR73 = {main_dev_in[99:0], 7'h49};
  ZLL_Main_dev2  instR73 (zll_main_dev2_inR73[106:7], zll_main_dev2_inR73[6:0], zll_main_dev2_outR73);
  assign zll_main_dev2_inR74 = {main_dev_in[99:0], 7'h4a};
  ZLL_Main_dev2  instR74 (zll_main_dev2_inR74[106:7], zll_main_dev2_inR74[6:0], zll_main_dev2_outR74);
  assign zll_main_dev2_inR75 = {main_dev_in[99:0], 7'h4b};
  ZLL_Main_dev2  instR75 (zll_main_dev2_inR75[106:7], zll_main_dev2_inR75[6:0], zll_main_dev2_outR75);
  assign zll_main_dev2_inR76 = {main_dev_in[99:0], 7'h4c};
  ZLL_Main_dev2  instR76 (zll_main_dev2_inR76[106:7], zll_main_dev2_inR76[6:0], zll_main_dev2_outR76);
  assign zll_main_dev2_inR77 = {main_dev_in[99:0], 7'h4d};
  ZLL_Main_dev2  instR77 (zll_main_dev2_inR77[106:7], zll_main_dev2_inR77[6:0], zll_main_dev2_outR77);
  assign zll_main_dev2_inR78 = {main_dev_in[99:0], 7'h4e};
  ZLL_Main_dev2  instR78 (zll_main_dev2_inR78[106:7], zll_main_dev2_inR78[6:0], zll_main_dev2_outR78);
  assign zll_main_dev2_inR79 = {main_dev_in[99:0], 7'h4f};
  ZLL_Main_dev2  instR79 (zll_main_dev2_inR79[106:7], zll_main_dev2_inR79[6:0], zll_main_dev2_outR79);
  assign zll_main_dev2_inR80 = {main_dev_in[99:0], 7'h50};
  ZLL_Main_dev2  instR80 (zll_main_dev2_inR80[106:7], zll_main_dev2_inR80[6:0], zll_main_dev2_outR80);
  assign zll_main_dev2_inR81 = {main_dev_in[99:0], 7'h51};
  ZLL_Main_dev2  instR81 (zll_main_dev2_inR81[106:7], zll_main_dev2_inR81[6:0], zll_main_dev2_outR81);
  assign zll_main_dev2_inR82 = {main_dev_in[99:0], 7'h52};
  ZLL_Main_dev2  instR82 (zll_main_dev2_inR82[106:7], zll_main_dev2_inR82[6:0], zll_main_dev2_outR82);
  assign zll_main_dev2_inR83 = {main_dev_in[99:0], 7'h53};
  ZLL_Main_dev2  instR83 (zll_main_dev2_inR83[106:7], zll_main_dev2_inR83[6:0], zll_main_dev2_outR83);
  assign zll_main_dev2_inR84 = {main_dev_in[99:0], 7'h54};
  ZLL_Main_dev2  instR84 (zll_main_dev2_inR84[106:7], zll_main_dev2_inR84[6:0], zll_main_dev2_outR84);
  assign zll_main_dev2_inR85 = {main_dev_in[99:0], 7'h55};
  ZLL_Main_dev2  instR85 (zll_main_dev2_inR85[106:7], zll_main_dev2_inR85[6:0], zll_main_dev2_outR85);
  assign zll_main_dev2_inR86 = {main_dev_in[99:0], 7'h56};
  ZLL_Main_dev2  instR86 (zll_main_dev2_inR86[106:7], zll_main_dev2_inR86[6:0], zll_main_dev2_outR86);
  assign zll_main_dev2_inR87 = {main_dev_in[99:0], 7'h57};
  ZLL_Main_dev2  instR87 (zll_main_dev2_inR87[106:7], zll_main_dev2_inR87[6:0], zll_main_dev2_outR87);
  assign zll_main_dev2_inR88 = {main_dev_in[99:0], 7'h58};
  ZLL_Main_dev2  instR88 (zll_main_dev2_inR88[106:7], zll_main_dev2_inR88[6:0], zll_main_dev2_outR88);
  assign zll_main_dev2_inR89 = {main_dev_in[99:0], 7'h59};
  ZLL_Main_dev2  instR89 (zll_main_dev2_inR89[106:7], zll_main_dev2_inR89[6:0], zll_main_dev2_outR89);
  assign zll_main_dev2_inR90 = {main_dev_in[99:0], 7'h5a};
  ZLL_Main_dev2  instR90 (zll_main_dev2_inR90[106:7], zll_main_dev2_inR90[6:0], zll_main_dev2_outR90);
  assign zll_main_dev2_inR91 = {main_dev_in[99:0], 7'h5b};
  ZLL_Main_dev2  instR91 (zll_main_dev2_inR91[106:7], zll_main_dev2_inR91[6:0], zll_main_dev2_outR91);
  assign zll_main_dev2_inR92 = {main_dev_in[99:0], 7'h5c};
  ZLL_Main_dev2  instR92 (zll_main_dev2_inR92[106:7], zll_main_dev2_inR92[6:0], zll_main_dev2_outR92);
  assign zll_main_dev2_inR93 = {main_dev_in[99:0], 7'h5d};
  ZLL_Main_dev2  instR93 (zll_main_dev2_inR93[106:7], zll_main_dev2_inR93[6:0], zll_main_dev2_outR93);
  assign zll_main_dev2_inR94 = {main_dev_in[99:0], 7'h5e};
  ZLL_Main_dev2  instR94 (zll_main_dev2_inR94[106:7], zll_main_dev2_inR94[6:0], zll_main_dev2_outR94);
  assign zll_main_dev2_inR95 = {main_dev_in[99:0], 7'h5f};
  ZLL_Main_dev2  instR95 (zll_main_dev2_inR95[106:7], zll_main_dev2_inR95[6:0], zll_main_dev2_outR95);
  assign zll_main_dev2_inR96 = {main_dev_in[99:0], 7'h60};
  ZLL_Main_dev2  instR96 (zll_main_dev2_inR96[106:7], zll_main_dev2_inR96[6:0], zll_main_dev2_outR96);
  assign zll_main_dev2_inR97 = {main_dev_in[99:0], 7'h61};
  ZLL_Main_dev2  instR97 (zll_main_dev2_inR97[106:7], zll_main_dev2_inR97[6:0], zll_main_dev2_outR97);
  assign zll_main_dev2_inR98 = {main_dev_in[99:0], 7'h62};
  ZLL_Main_dev2  instR98 (zll_main_dev2_inR98[106:7], zll_main_dev2_inR98[6:0], zll_main_dev2_outR98);
  assign zll_main_dev2_inR99 = {main_dev_in[99:0], 7'h63};
  ZLL_Main_dev2  instR99 (zll_main_dev2_inR99[106:7], zll_main_dev2_inR99[6:0], zll_main_dev2_outR99);
  assign zll_main_dev5_in = {main_dev_in[99:0], 7'h00};
  ZLL_Main_dev5  instR100 (zll_main_dev5_in[106:7], zll_main_dev5_in[6:0], zll_main_dev5_out);
  assign zll_main_dev5_inR1 = {main_dev_in[99:0], 7'h01};
  ZLL_Main_dev5  instR101 (zll_main_dev5_inR1[106:7], zll_main_dev5_inR1[6:0], zll_main_dev5_outR1);
  assign zll_main_dev5_inR2 = {main_dev_in[99:0], 7'h02};
  ZLL_Main_dev5  instR102 (zll_main_dev5_inR2[106:7], zll_main_dev5_inR2[6:0], zll_main_dev5_outR2);
  assign zll_main_dev5_inR3 = {main_dev_in[99:0], 7'h03};
  ZLL_Main_dev5  instR103 (zll_main_dev5_inR3[106:7], zll_main_dev5_inR3[6:0], zll_main_dev5_outR3);
  assign zll_main_dev5_inR4 = {main_dev_in[99:0], 7'h04};
  ZLL_Main_dev5  instR104 (zll_main_dev5_inR4[106:7], zll_main_dev5_inR4[6:0], zll_main_dev5_outR4);
  assign zll_main_dev5_inR5 = {main_dev_in[99:0], 7'h05};
  ZLL_Main_dev5  instR105 (zll_main_dev5_inR5[106:7], zll_main_dev5_inR5[6:0], zll_main_dev5_outR5);
  assign zll_main_dev5_inR6 = {main_dev_in[99:0], 7'h06};
  ZLL_Main_dev5  instR106 (zll_main_dev5_inR6[106:7], zll_main_dev5_inR6[6:0], zll_main_dev5_outR6);
  assign zll_main_dev5_inR7 = {main_dev_in[99:0], 7'h07};
  ZLL_Main_dev5  instR107 (zll_main_dev5_inR7[106:7], zll_main_dev5_inR7[6:0], zll_main_dev5_outR7);
  assign zll_main_dev5_inR8 = {main_dev_in[99:0], 7'h08};
  ZLL_Main_dev5  instR108 (zll_main_dev5_inR8[106:7], zll_main_dev5_inR8[6:0], zll_main_dev5_outR8);
  assign zll_main_dev5_inR9 = {main_dev_in[99:0], 7'h09};
  ZLL_Main_dev5  instR109 (zll_main_dev5_inR9[106:7], zll_main_dev5_inR9[6:0], zll_main_dev5_outR9);
  assign zll_main_dev5_inR10 = {main_dev_in[99:0], 7'h0a};
  ZLL_Main_dev5  instR110 (zll_main_dev5_inR10[106:7], zll_main_dev5_inR10[6:0], zll_main_dev5_outR10);
  assign zll_main_dev5_inR11 = {main_dev_in[99:0], 7'h0b};
  ZLL_Main_dev5  instR111 (zll_main_dev5_inR11[106:7], zll_main_dev5_inR11[6:0], zll_main_dev5_outR11);
  assign zll_main_dev5_inR12 = {main_dev_in[99:0], 7'h0c};
  ZLL_Main_dev5  instR112 (zll_main_dev5_inR12[106:7], zll_main_dev5_inR12[6:0], zll_main_dev5_outR12);
  assign zll_main_dev5_inR13 = {main_dev_in[99:0], 7'h0d};
  ZLL_Main_dev5  instR113 (zll_main_dev5_inR13[106:7], zll_main_dev5_inR13[6:0], zll_main_dev5_outR13);
  assign zll_main_dev5_inR14 = {main_dev_in[99:0], 7'h0e};
  ZLL_Main_dev5  instR114 (zll_main_dev5_inR14[106:7], zll_main_dev5_inR14[6:0], zll_main_dev5_outR14);
  assign zll_main_dev5_inR15 = {main_dev_in[99:0], 7'h0f};
  ZLL_Main_dev5  instR115 (zll_main_dev5_inR15[106:7], zll_main_dev5_inR15[6:0], zll_main_dev5_outR15);
  assign zll_main_dev5_inR16 = {main_dev_in[99:0], 7'h10};
  ZLL_Main_dev5  instR116 (zll_main_dev5_inR16[106:7], zll_main_dev5_inR16[6:0], zll_main_dev5_outR16);
  assign zll_main_dev5_inR17 = {main_dev_in[99:0], 7'h11};
  ZLL_Main_dev5  instR117 (zll_main_dev5_inR17[106:7], zll_main_dev5_inR17[6:0], zll_main_dev5_outR17);
  assign zll_main_dev5_inR18 = {main_dev_in[99:0], 7'h12};
  ZLL_Main_dev5  instR118 (zll_main_dev5_inR18[106:7], zll_main_dev5_inR18[6:0], zll_main_dev5_outR18);
  assign zll_main_dev5_inR19 = {main_dev_in[99:0], 7'h13};
  ZLL_Main_dev5  instR119 (zll_main_dev5_inR19[106:7], zll_main_dev5_inR19[6:0], zll_main_dev5_outR19);
  assign zll_main_dev5_inR20 = {main_dev_in[99:0], 7'h14};
  ZLL_Main_dev5  instR120 (zll_main_dev5_inR20[106:7], zll_main_dev5_inR20[6:0], zll_main_dev5_outR20);
  assign zll_main_dev5_inR21 = {main_dev_in[99:0], 7'h15};
  ZLL_Main_dev5  instR121 (zll_main_dev5_inR21[106:7], zll_main_dev5_inR21[6:0], zll_main_dev5_outR21);
  assign zll_main_dev5_inR22 = {main_dev_in[99:0], 7'h16};
  ZLL_Main_dev5  instR122 (zll_main_dev5_inR22[106:7], zll_main_dev5_inR22[6:0], zll_main_dev5_outR22);
  assign zll_main_dev5_inR23 = {main_dev_in[99:0], 7'h17};
  ZLL_Main_dev5  instR123 (zll_main_dev5_inR23[106:7], zll_main_dev5_inR23[6:0], zll_main_dev5_outR23);
  assign zll_main_dev5_inR24 = {main_dev_in[99:0], 7'h18};
  ZLL_Main_dev5  instR124 (zll_main_dev5_inR24[106:7], zll_main_dev5_inR24[6:0], zll_main_dev5_outR24);
  assign zll_main_dev5_inR25 = {main_dev_in[99:0], 7'h19};
  ZLL_Main_dev5  instR125 (zll_main_dev5_inR25[106:7], zll_main_dev5_inR25[6:0], zll_main_dev5_outR25);
  assign zll_main_dev5_inR26 = {main_dev_in[99:0], 7'h1a};
  ZLL_Main_dev5  instR126 (zll_main_dev5_inR26[106:7], zll_main_dev5_inR26[6:0], zll_main_dev5_outR26);
  assign zll_main_dev5_inR27 = {main_dev_in[99:0], 7'h1b};
  ZLL_Main_dev5  instR127 (zll_main_dev5_inR27[106:7], zll_main_dev5_inR27[6:0], zll_main_dev5_outR27);
  assign zll_main_dev5_inR28 = {main_dev_in[99:0], 7'h1c};
  ZLL_Main_dev5  instR128 (zll_main_dev5_inR28[106:7], zll_main_dev5_inR28[6:0], zll_main_dev5_outR28);
  assign zll_main_dev5_inR29 = {main_dev_in[99:0], 7'h1d};
  ZLL_Main_dev5  instR129 (zll_main_dev5_inR29[106:7], zll_main_dev5_inR29[6:0], zll_main_dev5_outR29);
  assign zll_main_dev5_inR30 = {main_dev_in[99:0], 7'h1e};
  ZLL_Main_dev5  instR130 (zll_main_dev5_inR30[106:7], zll_main_dev5_inR30[6:0], zll_main_dev5_outR30);
  assign zll_main_dev5_inR31 = {main_dev_in[99:0], 7'h1f};
  ZLL_Main_dev5  instR131 (zll_main_dev5_inR31[106:7], zll_main_dev5_inR31[6:0], zll_main_dev5_outR31);
  assign zll_main_dev5_inR32 = {main_dev_in[99:0], 7'h20};
  ZLL_Main_dev5  instR132 (zll_main_dev5_inR32[106:7], zll_main_dev5_inR32[6:0], zll_main_dev5_outR32);
  assign zll_main_dev5_inR33 = {main_dev_in[99:0], 7'h21};
  ZLL_Main_dev5  instR133 (zll_main_dev5_inR33[106:7], zll_main_dev5_inR33[6:0], zll_main_dev5_outR33);
  assign zll_main_dev5_inR34 = {main_dev_in[99:0], 7'h22};
  ZLL_Main_dev5  instR134 (zll_main_dev5_inR34[106:7], zll_main_dev5_inR34[6:0], zll_main_dev5_outR34);
  assign zll_main_dev5_inR35 = {main_dev_in[99:0], 7'h23};
  ZLL_Main_dev5  instR135 (zll_main_dev5_inR35[106:7], zll_main_dev5_inR35[6:0], zll_main_dev5_outR35);
  assign zll_main_dev5_inR36 = {main_dev_in[99:0], 7'h24};
  ZLL_Main_dev5  instR136 (zll_main_dev5_inR36[106:7], zll_main_dev5_inR36[6:0], zll_main_dev5_outR36);
  assign zll_main_dev5_inR37 = {main_dev_in[99:0], 7'h25};
  ZLL_Main_dev5  instR137 (zll_main_dev5_inR37[106:7], zll_main_dev5_inR37[6:0], zll_main_dev5_outR37);
  assign zll_main_dev5_inR38 = {main_dev_in[99:0], 7'h26};
  ZLL_Main_dev5  instR138 (zll_main_dev5_inR38[106:7], zll_main_dev5_inR38[6:0], zll_main_dev5_outR38);
  assign zll_main_dev5_inR39 = {main_dev_in[99:0], 7'h27};
  ZLL_Main_dev5  instR139 (zll_main_dev5_inR39[106:7], zll_main_dev5_inR39[6:0], zll_main_dev5_outR39);
  assign zll_main_dev5_inR40 = {main_dev_in[99:0], 7'h28};
  ZLL_Main_dev5  instR140 (zll_main_dev5_inR40[106:7], zll_main_dev5_inR40[6:0], zll_main_dev5_outR40);
  assign zll_main_dev5_inR41 = {main_dev_in[99:0], 7'h29};
  ZLL_Main_dev5  instR141 (zll_main_dev5_inR41[106:7], zll_main_dev5_inR41[6:0], zll_main_dev5_outR41);
  assign zll_main_dev5_inR42 = {main_dev_in[99:0], 7'h2a};
  ZLL_Main_dev5  instR142 (zll_main_dev5_inR42[106:7], zll_main_dev5_inR42[6:0], zll_main_dev5_outR42);
  assign zll_main_dev5_inR43 = {main_dev_in[99:0], 7'h2b};
  ZLL_Main_dev5  instR143 (zll_main_dev5_inR43[106:7], zll_main_dev5_inR43[6:0], zll_main_dev5_outR43);
  assign zll_main_dev5_inR44 = {main_dev_in[99:0], 7'h2c};
  ZLL_Main_dev5  instR144 (zll_main_dev5_inR44[106:7], zll_main_dev5_inR44[6:0], zll_main_dev5_outR44);
  assign zll_main_dev5_inR45 = {main_dev_in[99:0], 7'h2d};
  ZLL_Main_dev5  instR145 (zll_main_dev5_inR45[106:7], zll_main_dev5_inR45[6:0], zll_main_dev5_outR45);
  assign zll_main_dev5_inR46 = {main_dev_in[99:0], 7'h2e};
  ZLL_Main_dev5  instR146 (zll_main_dev5_inR46[106:7], zll_main_dev5_inR46[6:0], zll_main_dev5_outR46);
  assign zll_main_dev5_inR47 = {main_dev_in[99:0], 7'h2f};
  ZLL_Main_dev5  instR147 (zll_main_dev5_inR47[106:7], zll_main_dev5_inR47[6:0], zll_main_dev5_outR47);
  assign zll_main_dev5_inR48 = {main_dev_in[99:0], 7'h30};
  ZLL_Main_dev5  instR148 (zll_main_dev5_inR48[106:7], zll_main_dev5_inR48[6:0], zll_main_dev5_outR48);
  assign zll_main_dev5_inR49 = {main_dev_in[99:0], 7'h31};
  ZLL_Main_dev5  instR149 (zll_main_dev5_inR49[106:7], zll_main_dev5_inR49[6:0], zll_main_dev5_outR49);
  assign zll_main_dev5_inR50 = {main_dev_in[99:0], 7'h32};
  ZLL_Main_dev5  instR150 (zll_main_dev5_inR50[106:7], zll_main_dev5_inR50[6:0], zll_main_dev5_outR50);
  assign zll_main_dev5_inR51 = {main_dev_in[99:0], 7'h33};
  ZLL_Main_dev5  instR151 (zll_main_dev5_inR51[106:7], zll_main_dev5_inR51[6:0], zll_main_dev5_outR51);
  assign zll_main_dev5_inR52 = {main_dev_in[99:0], 7'h34};
  ZLL_Main_dev5  instR152 (zll_main_dev5_inR52[106:7], zll_main_dev5_inR52[6:0], zll_main_dev5_outR52);
  assign zll_main_dev5_inR53 = {main_dev_in[99:0], 7'h35};
  ZLL_Main_dev5  instR153 (zll_main_dev5_inR53[106:7], zll_main_dev5_inR53[6:0], zll_main_dev5_outR53);
  assign zll_main_dev5_inR54 = {main_dev_in[99:0], 7'h36};
  ZLL_Main_dev5  instR154 (zll_main_dev5_inR54[106:7], zll_main_dev5_inR54[6:0], zll_main_dev5_outR54);
  assign zll_main_dev5_inR55 = {main_dev_in[99:0], 7'h37};
  ZLL_Main_dev5  instR155 (zll_main_dev5_inR55[106:7], zll_main_dev5_inR55[6:0], zll_main_dev5_outR55);
  assign zll_main_dev5_inR56 = {main_dev_in[99:0], 7'h38};
  ZLL_Main_dev5  instR156 (zll_main_dev5_inR56[106:7], zll_main_dev5_inR56[6:0], zll_main_dev5_outR56);
  assign zll_main_dev5_inR57 = {main_dev_in[99:0], 7'h39};
  ZLL_Main_dev5  instR157 (zll_main_dev5_inR57[106:7], zll_main_dev5_inR57[6:0], zll_main_dev5_outR57);
  assign zll_main_dev5_inR58 = {main_dev_in[99:0], 7'h3a};
  ZLL_Main_dev5  instR158 (zll_main_dev5_inR58[106:7], zll_main_dev5_inR58[6:0], zll_main_dev5_outR58);
  assign zll_main_dev5_inR59 = {main_dev_in[99:0], 7'h3b};
  ZLL_Main_dev5  instR159 (zll_main_dev5_inR59[106:7], zll_main_dev5_inR59[6:0], zll_main_dev5_outR59);
  assign zll_main_dev5_inR60 = {main_dev_in[99:0], 7'h3c};
  ZLL_Main_dev5  instR160 (zll_main_dev5_inR60[106:7], zll_main_dev5_inR60[6:0], zll_main_dev5_outR60);
  assign zll_main_dev5_inR61 = {main_dev_in[99:0], 7'h3d};
  ZLL_Main_dev5  instR161 (zll_main_dev5_inR61[106:7], zll_main_dev5_inR61[6:0], zll_main_dev5_outR61);
  assign zll_main_dev5_inR62 = {main_dev_in[99:0], 7'h3e};
  ZLL_Main_dev5  instR162 (zll_main_dev5_inR62[106:7], zll_main_dev5_inR62[6:0], zll_main_dev5_outR62);
  assign zll_main_dev5_inR63 = {main_dev_in[99:0], 7'h3f};
  ZLL_Main_dev5  instR163 (zll_main_dev5_inR63[106:7], zll_main_dev5_inR63[6:0], zll_main_dev5_outR63);
  assign zll_main_dev5_inR64 = {main_dev_in[99:0], 7'h40};
  ZLL_Main_dev5  instR164 (zll_main_dev5_inR64[106:7], zll_main_dev5_inR64[6:0], zll_main_dev5_outR64);
  assign zll_main_dev5_inR65 = {main_dev_in[99:0], 7'h41};
  ZLL_Main_dev5  instR165 (zll_main_dev5_inR65[106:7], zll_main_dev5_inR65[6:0], zll_main_dev5_outR65);
  assign zll_main_dev5_inR66 = {main_dev_in[99:0], 7'h42};
  ZLL_Main_dev5  instR166 (zll_main_dev5_inR66[106:7], zll_main_dev5_inR66[6:0], zll_main_dev5_outR66);
  assign zll_main_dev5_inR67 = {main_dev_in[99:0], 7'h43};
  ZLL_Main_dev5  instR167 (zll_main_dev5_inR67[106:7], zll_main_dev5_inR67[6:0], zll_main_dev5_outR67);
  assign zll_main_dev5_inR68 = {main_dev_in[99:0], 7'h44};
  ZLL_Main_dev5  instR168 (zll_main_dev5_inR68[106:7], zll_main_dev5_inR68[6:0], zll_main_dev5_outR68);
  assign zll_main_dev5_inR69 = {main_dev_in[99:0], 7'h45};
  ZLL_Main_dev5  instR169 (zll_main_dev5_inR69[106:7], zll_main_dev5_inR69[6:0], zll_main_dev5_outR69);
  assign zll_main_dev5_inR70 = {main_dev_in[99:0], 7'h46};
  ZLL_Main_dev5  instR170 (zll_main_dev5_inR70[106:7], zll_main_dev5_inR70[6:0], zll_main_dev5_outR70);
  assign zll_main_dev5_inR71 = {main_dev_in[99:0], 7'h47};
  ZLL_Main_dev5  instR171 (zll_main_dev5_inR71[106:7], zll_main_dev5_inR71[6:0], zll_main_dev5_outR71);
  assign zll_main_dev5_inR72 = {main_dev_in[99:0], 7'h48};
  ZLL_Main_dev5  instR172 (zll_main_dev5_inR72[106:7], zll_main_dev5_inR72[6:0], zll_main_dev5_outR72);
  assign zll_main_dev5_inR73 = {main_dev_in[99:0], 7'h49};
  ZLL_Main_dev5  instR173 (zll_main_dev5_inR73[106:7], zll_main_dev5_inR73[6:0], zll_main_dev5_outR73);
  assign zll_main_dev5_inR74 = {main_dev_in[99:0], 7'h4a};
  ZLL_Main_dev5  instR174 (zll_main_dev5_inR74[106:7], zll_main_dev5_inR74[6:0], zll_main_dev5_outR74);
  assign zll_main_dev5_inR75 = {main_dev_in[99:0], 7'h4b};
  ZLL_Main_dev5  instR175 (zll_main_dev5_inR75[106:7], zll_main_dev5_inR75[6:0], zll_main_dev5_outR75);
  assign zll_main_dev5_inR76 = {main_dev_in[99:0], 7'h4c};
  ZLL_Main_dev5  instR176 (zll_main_dev5_inR76[106:7], zll_main_dev5_inR76[6:0], zll_main_dev5_outR76);
  assign zll_main_dev5_inR77 = {main_dev_in[99:0], 7'h4d};
  ZLL_Main_dev5  instR177 (zll_main_dev5_inR77[106:7], zll_main_dev5_inR77[6:0], zll_main_dev5_outR77);
  assign zll_main_dev5_inR78 = {main_dev_in[99:0], 7'h4e};
  ZLL_Main_dev5  instR178 (zll_main_dev5_inR78[106:7], zll_main_dev5_inR78[6:0], zll_main_dev5_outR78);
  assign zll_main_dev5_inR79 = {main_dev_in[99:0], 7'h4f};
  ZLL_Main_dev5  instR179 (zll_main_dev5_inR79[106:7], zll_main_dev5_inR79[6:0], zll_main_dev5_outR79);
  assign zll_main_dev5_inR80 = {main_dev_in[99:0], 7'h50};
  ZLL_Main_dev5  instR180 (zll_main_dev5_inR80[106:7], zll_main_dev5_inR80[6:0], zll_main_dev5_outR80);
  assign zll_main_dev5_inR81 = {main_dev_in[99:0], 7'h51};
  ZLL_Main_dev5  instR181 (zll_main_dev5_inR81[106:7], zll_main_dev5_inR81[6:0], zll_main_dev5_outR81);
  assign zll_main_dev5_inR82 = {main_dev_in[99:0], 7'h52};
  ZLL_Main_dev5  instR182 (zll_main_dev5_inR82[106:7], zll_main_dev5_inR82[6:0], zll_main_dev5_outR82);
  assign zll_main_dev5_inR83 = {main_dev_in[99:0], 7'h53};
  ZLL_Main_dev5  instR183 (zll_main_dev5_inR83[106:7], zll_main_dev5_inR83[6:0], zll_main_dev5_outR83);
  assign zll_main_dev5_inR84 = {main_dev_in[99:0], 7'h54};
  ZLL_Main_dev5  instR184 (zll_main_dev5_inR84[106:7], zll_main_dev5_inR84[6:0], zll_main_dev5_outR84);
  assign zll_main_dev5_inR85 = {main_dev_in[99:0], 7'h55};
  ZLL_Main_dev5  instR185 (zll_main_dev5_inR85[106:7], zll_main_dev5_inR85[6:0], zll_main_dev5_outR85);
  assign zll_main_dev5_inR86 = {main_dev_in[99:0], 7'h56};
  ZLL_Main_dev5  instR186 (zll_main_dev5_inR86[106:7], zll_main_dev5_inR86[6:0], zll_main_dev5_outR86);
  assign zll_main_dev5_inR87 = {main_dev_in[99:0], 7'h57};
  ZLL_Main_dev5  instR187 (zll_main_dev5_inR87[106:7], zll_main_dev5_inR87[6:0], zll_main_dev5_outR87);
  assign zll_main_dev5_inR88 = {main_dev_in[99:0], 7'h58};
  ZLL_Main_dev5  instR188 (zll_main_dev5_inR88[106:7], zll_main_dev5_inR88[6:0], zll_main_dev5_outR88);
  assign zll_main_dev5_inR89 = {main_dev_in[99:0], 7'h59};
  ZLL_Main_dev5  instR189 (zll_main_dev5_inR89[106:7], zll_main_dev5_inR89[6:0], zll_main_dev5_outR89);
  assign zll_main_dev5_inR90 = {main_dev_in[99:0], 7'h5a};
  ZLL_Main_dev5  instR190 (zll_main_dev5_inR90[106:7], zll_main_dev5_inR90[6:0], zll_main_dev5_outR90);
  assign zll_main_dev5_inR91 = {main_dev_in[99:0], 7'h5b};
  ZLL_Main_dev5  instR191 (zll_main_dev5_inR91[106:7], zll_main_dev5_inR91[6:0], zll_main_dev5_outR91);
  assign zll_main_dev5_inR92 = {main_dev_in[99:0], 7'h5c};
  ZLL_Main_dev5  instR192 (zll_main_dev5_inR92[106:7], zll_main_dev5_inR92[6:0], zll_main_dev5_outR92);
  assign zll_main_dev5_inR93 = {main_dev_in[99:0], 7'h5d};
  ZLL_Main_dev5  instR193 (zll_main_dev5_inR93[106:7], zll_main_dev5_inR93[6:0], zll_main_dev5_outR93);
  assign zll_main_dev5_inR94 = {main_dev_in[99:0], 7'h5e};
  ZLL_Main_dev5  instR194 (zll_main_dev5_inR94[106:7], zll_main_dev5_inR94[6:0], zll_main_dev5_outR94);
  assign zll_main_dev5_inR95 = {main_dev_in[99:0], 7'h5f};
  ZLL_Main_dev5  instR195 (zll_main_dev5_inR95[106:7], zll_main_dev5_inR95[6:0], zll_main_dev5_outR95);
  assign zll_main_dev5_inR96 = {main_dev_in[99:0], 7'h60};
  ZLL_Main_dev5  instR196 (zll_main_dev5_inR96[106:7], zll_main_dev5_inR96[6:0], zll_main_dev5_outR96);
  assign zll_main_dev5_inR97 = {main_dev_in[99:0], 7'h61};
  ZLL_Main_dev5  instR197 (zll_main_dev5_inR97[106:7], zll_main_dev5_inR97[6:0], zll_main_dev5_outR97);
  assign zll_main_dev5_inR98 = {main_dev_in[99:0], 7'h62};
  ZLL_Main_dev5  instR198 (zll_main_dev5_inR98[106:7], zll_main_dev5_inR98[6:0], zll_main_dev5_outR98);
  assign zll_main_dev5_inR99 = {main_dev_in[99:0], 7'h63};
  ZLL_Main_dev5  instR199 (zll_main_dev5_inR99[106:7], zll_main_dev5_inR99[6:0], zll_main_dev5_outR99);
  assign zll_main_dev8_in = {main_dev_in[99:0], 7'h00};
  ZLL_Main_dev8  instR200 (zll_main_dev8_in[106:7], zll_main_dev8_in[6:0], zll_main_dev8_out);
  assign zll_main_dev8_inR1 = {main_dev_in[99:0], 7'h01};
  ZLL_Main_dev8  instR201 (zll_main_dev8_inR1[106:7], zll_main_dev8_inR1[6:0], zll_main_dev8_outR1);
  assign zll_main_dev8_inR2 = {main_dev_in[99:0], 7'h02};
  ZLL_Main_dev8  instR202 (zll_main_dev8_inR2[106:7], zll_main_dev8_inR2[6:0], zll_main_dev8_outR2);
  assign zll_main_dev8_inR3 = {main_dev_in[99:0], 7'h03};
  ZLL_Main_dev8  instR203 (zll_main_dev8_inR3[106:7], zll_main_dev8_inR3[6:0], zll_main_dev8_outR3);
  assign zll_main_dev8_inR4 = {main_dev_in[99:0], 7'h04};
  ZLL_Main_dev8  instR204 (zll_main_dev8_inR4[106:7], zll_main_dev8_inR4[6:0], zll_main_dev8_outR4);
  assign zll_main_dev8_inR5 = {main_dev_in[99:0], 7'h05};
  ZLL_Main_dev8  instR205 (zll_main_dev8_inR5[106:7], zll_main_dev8_inR5[6:0], zll_main_dev8_outR5);
  assign zll_main_dev8_inR6 = {main_dev_in[99:0], 7'h06};
  ZLL_Main_dev8  instR206 (zll_main_dev8_inR6[106:7], zll_main_dev8_inR6[6:0], zll_main_dev8_outR6);
  assign zll_main_dev8_inR7 = {main_dev_in[99:0], 7'h07};
  ZLL_Main_dev8  instR207 (zll_main_dev8_inR7[106:7], zll_main_dev8_inR7[6:0], zll_main_dev8_outR7);
  assign zll_main_dev8_inR8 = {main_dev_in[99:0], 7'h08};
  ZLL_Main_dev8  instR208 (zll_main_dev8_inR8[106:7], zll_main_dev8_inR8[6:0], zll_main_dev8_outR8);
  assign zll_main_dev8_inR9 = {main_dev_in[99:0], 7'h09};
  ZLL_Main_dev8  instR209 (zll_main_dev8_inR9[106:7], zll_main_dev8_inR9[6:0], zll_main_dev8_outR9);
  assign zll_main_dev8_inR10 = {main_dev_in[99:0], 7'h0a};
  ZLL_Main_dev8  instR210 (zll_main_dev8_inR10[106:7], zll_main_dev8_inR10[6:0], zll_main_dev8_outR10);
  assign zll_main_dev8_inR11 = {main_dev_in[99:0], 7'h0b};
  ZLL_Main_dev8  instR211 (zll_main_dev8_inR11[106:7], zll_main_dev8_inR11[6:0], zll_main_dev8_outR11);
  assign zll_main_dev8_inR12 = {main_dev_in[99:0], 7'h0c};
  ZLL_Main_dev8  instR212 (zll_main_dev8_inR12[106:7], zll_main_dev8_inR12[6:0], zll_main_dev8_outR12);
  assign zll_main_dev8_inR13 = {main_dev_in[99:0], 7'h0d};
  ZLL_Main_dev8  instR213 (zll_main_dev8_inR13[106:7], zll_main_dev8_inR13[6:0], zll_main_dev8_outR13);
  assign zll_main_dev8_inR14 = {main_dev_in[99:0], 7'h0e};
  ZLL_Main_dev8  instR214 (zll_main_dev8_inR14[106:7], zll_main_dev8_inR14[6:0], zll_main_dev8_outR14);
  assign zll_main_dev8_inR15 = {main_dev_in[99:0], 7'h0f};
  ZLL_Main_dev8  instR215 (zll_main_dev8_inR15[106:7], zll_main_dev8_inR15[6:0], zll_main_dev8_outR15);
  assign zll_main_dev8_inR16 = {main_dev_in[99:0], 7'h10};
  ZLL_Main_dev8  instR216 (zll_main_dev8_inR16[106:7], zll_main_dev8_inR16[6:0], zll_main_dev8_outR16);
  assign zll_main_dev8_inR17 = {main_dev_in[99:0], 7'h11};
  ZLL_Main_dev8  instR217 (zll_main_dev8_inR17[106:7], zll_main_dev8_inR17[6:0], zll_main_dev8_outR17);
  assign zll_main_dev8_inR18 = {main_dev_in[99:0], 7'h12};
  ZLL_Main_dev8  instR218 (zll_main_dev8_inR18[106:7], zll_main_dev8_inR18[6:0], zll_main_dev8_outR18);
  assign zll_main_dev8_inR19 = {main_dev_in[99:0], 7'h13};
  ZLL_Main_dev8  instR219 (zll_main_dev8_inR19[106:7], zll_main_dev8_inR19[6:0], zll_main_dev8_outR19);
  assign zll_main_dev8_inR20 = {main_dev_in[99:0], 7'h14};
  ZLL_Main_dev8  instR220 (zll_main_dev8_inR20[106:7], zll_main_dev8_inR20[6:0], zll_main_dev8_outR20);
  assign zll_main_dev8_inR21 = {main_dev_in[99:0], 7'h15};
  ZLL_Main_dev8  instR221 (zll_main_dev8_inR21[106:7], zll_main_dev8_inR21[6:0], zll_main_dev8_outR21);
  assign zll_main_dev8_inR22 = {main_dev_in[99:0], 7'h16};
  ZLL_Main_dev8  instR222 (zll_main_dev8_inR22[106:7], zll_main_dev8_inR22[6:0], zll_main_dev8_outR22);
  assign zll_main_dev8_inR23 = {main_dev_in[99:0], 7'h17};
  ZLL_Main_dev8  instR223 (zll_main_dev8_inR23[106:7], zll_main_dev8_inR23[6:0], zll_main_dev8_outR23);
  assign zll_main_dev8_inR24 = {main_dev_in[99:0], 7'h18};
  ZLL_Main_dev8  instR224 (zll_main_dev8_inR24[106:7], zll_main_dev8_inR24[6:0], zll_main_dev8_outR24);
  assign zll_main_dev8_inR25 = {main_dev_in[99:0], 7'h19};
  ZLL_Main_dev8  instR225 (zll_main_dev8_inR25[106:7], zll_main_dev8_inR25[6:0], zll_main_dev8_outR25);
  assign zll_main_dev8_inR26 = {main_dev_in[99:0], 7'h1a};
  ZLL_Main_dev8  instR226 (zll_main_dev8_inR26[106:7], zll_main_dev8_inR26[6:0], zll_main_dev8_outR26);
  assign zll_main_dev8_inR27 = {main_dev_in[99:0], 7'h1b};
  ZLL_Main_dev8  instR227 (zll_main_dev8_inR27[106:7], zll_main_dev8_inR27[6:0], zll_main_dev8_outR27);
  assign zll_main_dev8_inR28 = {main_dev_in[99:0], 7'h1c};
  ZLL_Main_dev8  instR228 (zll_main_dev8_inR28[106:7], zll_main_dev8_inR28[6:0], zll_main_dev8_outR28);
  assign zll_main_dev8_inR29 = {main_dev_in[99:0], 7'h1d};
  ZLL_Main_dev8  instR229 (zll_main_dev8_inR29[106:7], zll_main_dev8_inR29[6:0], zll_main_dev8_outR29);
  assign zll_main_dev8_inR30 = {main_dev_in[99:0], 7'h1e};
  ZLL_Main_dev8  instR230 (zll_main_dev8_inR30[106:7], zll_main_dev8_inR30[6:0], zll_main_dev8_outR30);
  assign zll_main_dev8_inR31 = {main_dev_in[99:0], 7'h1f};
  ZLL_Main_dev8  instR231 (zll_main_dev8_inR31[106:7], zll_main_dev8_inR31[6:0], zll_main_dev8_outR31);
  assign zll_main_dev8_inR32 = {main_dev_in[99:0], 7'h20};
  ZLL_Main_dev8  instR232 (zll_main_dev8_inR32[106:7], zll_main_dev8_inR32[6:0], zll_main_dev8_outR32);
  assign zll_main_dev8_inR33 = {main_dev_in[99:0], 7'h21};
  ZLL_Main_dev8  instR233 (zll_main_dev8_inR33[106:7], zll_main_dev8_inR33[6:0], zll_main_dev8_outR33);
  assign zll_main_dev8_inR34 = {main_dev_in[99:0], 7'h22};
  ZLL_Main_dev8  instR234 (zll_main_dev8_inR34[106:7], zll_main_dev8_inR34[6:0], zll_main_dev8_outR34);
  assign zll_main_dev8_inR35 = {main_dev_in[99:0], 7'h23};
  ZLL_Main_dev8  instR235 (zll_main_dev8_inR35[106:7], zll_main_dev8_inR35[6:0], zll_main_dev8_outR35);
  assign zll_main_dev8_inR36 = {main_dev_in[99:0], 7'h24};
  ZLL_Main_dev8  instR236 (zll_main_dev8_inR36[106:7], zll_main_dev8_inR36[6:0], zll_main_dev8_outR36);
  assign zll_main_dev8_inR37 = {main_dev_in[99:0], 7'h25};
  ZLL_Main_dev8  instR237 (zll_main_dev8_inR37[106:7], zll_main_dev8_inR37[6:0], zll_main_dev8_outR37);
  assign zll_main_dev8_inR38 = {main_dev_in[99:0], 7'h26};
  ZLL_Main_dev8  instR238 (zll_main_dev8_inR38[106:7], zll_main_dev8_inR38[6:0], zll_main_dev8_outR38);
  assign zll_main_dev8_inR39 = {main_dev_in[99:0], 7'h27};
  ZLL_Main_dev8  instR239 (zll_main_dev8_inR39[106:7], zll_main_dev8_inR39[6:0], zll_main_dev8_outR39);
  assign zll_main_dev8_inR40 = {main_dev_in[99:0], 7'h28};
  ZLL_Main_dev8  instR240 (zll_main_dev8_inR40[106:7], zll_main_dev8_inR40[6:0], zll_main_dev8_outR40);
  assign zll_main_dev8_inR41 = {main_dev_in[99:0], 7'h29};
  ZLL_Main_dev8  instR241 (zll_main_dev8_inR41[106:7], zll_main_dev8_inR41[6:0], zll_main_dev8_outR41);
  assign zll_main_dev8_inR42 = {main_dev_in[99:0], 7'h2a};
  ZLL_Main_dev8  instR242 (zll_main_dev8_inR42[106:7], zll_main_dev8_inR42[6:0], zll_main_dev8_outR42);
  assign zll_main_dev8_inR43 = {main_dev_in[99:0], 7'h2b};
  ZLL_Main_dev8  instR243 (zll_main_dev8_inR43[106:7], zll_main_dev8_inR43[6:0], zll_main_dev8_outR43);
  assign zll_main_dev8_inR44 = {main_dev_in[99:0], 7'h2c};
  ZLL_Main_dev8  instR244 (zll_main_dev8_inR44[106:7], zll_main_dev8_inR44[6:0], zll_main_dev8_outR44);
  assign zll_main_dev8_inR45 = {main_dev_in[99:0], 7'h2d};
  ZLL_Main_dev8  instR245 (zll_main_dev8_inR45[106:7], zll_main_dev8_inR45[6:0], zll_main_dev8_outR45);
  assign zll_main_dev8_inR46 = {main_dev_in[99:0], 7'h2e};
  ZLL_Main_dev8  instR246 (zll_main_dev8_inR46[106:7], zll_main_dev8_inR46[6:0], zll_main_dev8_outR46);
  assign zll_main_dev8_inR47 = {main_dev_in[99:0], 7'h2f};
  ZLL_Main_dev8  instR247 (zll_main_dev8_inR47[106:7], zll_main_dev8_inR47[6:0], zll_main_dev8_outR47);
  assign zll_main_dev8_inR48 = {main_dev_in[99:0], 7'h30};
  ZLL_Main_dev8  instR248 (zll_main_dev8_inR48[106:7], zll_main_dev8_inR48[6:0], zll_main_dev8_outR48);
  assign zll_main_dev8_inR49 = {main_dev_in[99:0], 7'h31};
  ZLL_Main_dev8  instR249 (zll_main_dev8_inR49[106:7], zll_main_dev8_inR49[6:0], zll_main_dev8_outR49);
  assign zll_main_dev8_inR50 = {main_dev_in[99:0], 7'h32};
  ZLL_Main_dev8  instR250 (zll_main_dev8_inR50[106:7], zll_main_dev8_inR50[6:0], zll_main_dev8_outR50);
  assign zll_main_dev8_inR51 = {main_dev_in[99:0], 7'h33};
  ZLL_Main_dev8  instR251 (zll_main_dev8_inR51[106:7], zll_main_dev8_inR51[6:0], zll_main_dev8_outR51);
  assign zll_main_dev8_inR52 = {main_dev_in[99:0], 7'h34};
  ZLL_Main_dev8  instR252 (zll_main_dev8_inR52[106:7], zll_main_dev8_inR52[6:0], zll_main_dev8_outR52);
  assign zll_main_dev8_inR53 = {main_dev_in[99:0], 7'h35};
  ZLL_Main_dev8  instR253 (zll_main_dev8_inR53[106:7], zll_main_dev8_inR53[6:0], zll_main_dev8_outR53);
  assign zll_main_dev8_inR54 = {main_dev_in[99:0], 7'h36};
  ZLL_Main_dev8  instR254 (zll_main_dev8_inR54[106:7], zll_main_dev8_inR54[6:0], zll_main_dev8_outR54);
  assign zll_main_dev8_inR55 = {main_dev_in[99:0], 7'h37};
  ZLL_Main_dev8  instR255 (zll_main_dev8_inR55[106:7], zll_main_dev8_inR55[6:0], zll_main_dev8_outR55);
  assign zll_main_dev8_inR56 = {main_dev_in[99:0], 7'h38};
  ZLL_Main_dev8  instR256 (zll_main_dev8_inR56[106:7], zll_main_dev8_inR56[6:0], zll_main_dev8_outR56);
  assign zll_main_dev8_inR57 = {main_dev_in[99:0], 7'h39};
  ZLL_Main_dev8  instR257 (zll_main_dev8_inR57[106:7], zll_main_dev8_inR57[6:0], zll_main_dev8_outR57);
  assign zll_main_dev8_inR58 = {main_dev_in[99:0], 7'h3a};
  ZLL_Main_dev8  instR258 (zll_main_dev8_inR58[106:7], zll_main_dev8_inR58[6:0], zll_main_dev8_outR58);
  assign zll_main_dev8_inR59 = {main_dev_in[99:0], 7'h3b};
  ZLL_Main_dev8  instR259 (zll_main_dev8_inR59[106:7], zll_main_dev8_inR59[6:0], zll_main_dev8_outR59);
  assign zll_main_dev8_inR60 = {main_dev_in[99:0], 7'h3c};
  ZLL_Main_dev8  instR260 (zll_main_dev8_inR60[106:7], zll_main_dev8_inR60[6:0], zll_main_dev8_outR60);
  assign zll_main_dev8_inR61 = {main_dev_in[99:0], 7'h3d};
  ZLL_Main_dev8  instR261 (zll_main_dev8_inR61[106:7], zll_main_dev8_inR61[6:0], zll_main_dev8_outR61);
  assign zll_main_dev8_inR62 = {main_dev_in[99:0], 7'h3e};
  ZLL_Main_dev8  instR262 (zll_main_dev8_inR62[106:7], zll_main_dev8_inR62[6:0], zll_main_dev8_outR62);
  assign zll_main_dev8_inR63 = {main_dev_in[99:0], 7'h3f};
  ZLL_Main_dev8  instR263 (zll_main_dev8_inR63[106:7], zll_main_dev8_inR63[6:0], zll_main_dev8_outR63);
  assign zll_main_dev8_inR64 = {main_dev_in[99:0], 7'h40};
  ZLL_Main_dev8  instR264 (zll_main_dev8_inR64[106:7], zll_main_dev8_inR64[6:0], zll_main_dev8_outR64);
  assign zll_main_dev8_inR65 = {main_dev_in[99:0], 7'h41};
  ZLL_Main_dev8  instR265 (zll_main_dev8_inR65[106:7], zll_main_dev8_inR65[6:0], zll_main_dev8_outR65);
  assign zll_main_dev8_inR66 = {main_dev_in[99:0], 7'h42};
  ZLL_Main_dev8  instR266 (zll_main_dev8_inR66[106:7], zll_main_dev8_inR66[6:0], zll_main_dev8_outR66);
  assign zll_main_dev8_inR67 = {main_dev_in[99:0], 7'h43};
  ZLL_Main_dev8  instR267 (zll_main_dev8_inR67[106:7], zll_main_dev8_inR67[6:0], zll_main_dev8_outR67);
  assign zll_main_dev8_inR68 = {main_dev_in[99:0], 7'h44};
  ZLL_Main_dev8  instR268 (zll_main_dev8_inR68[106:7], zll_main_dev8_inR68[6:0], zll_main_dev8_outR68);
  assign zll_main_dev8_inR69 = {main_dev_in[99:0], 7'h45};
  ZLL_Main_dev8  instR269 (zll_main_dev8_inR69[106:7], zll_main_dev8_inR69[6:0], zll_main_dev8_outR69);
  assign zll_main_dev8_inR70 = {main_dev_in[99:0], 7'h46};
  ZLL_Main_dev8  instR270 (zll_main_dev8_inR70[106:7], zll_main_dev8_inR70[6:0], zll_main_dev8_outR70);
  assign zll_main_dev8_inR71 = {main_dev_in[99:0], 7'h47};
  ZLL_Main_dev8  instR271 (zll_main_dev8_inR71[106:7], zll_main_dev8_inR71[6:0], zll_main_dev8_outR71);
  assign zll_main_dev8_inR72 = {main_dev_in[99:0], 7'h48};
  ZLL_Main_dev8  instR272 (zll_main_dev8_inR72[106:7], zll_main_dev8_inR72[6:0], zll_main_dev8_outR72);
  assign zll_main_dev8_inR73 = {main_dev_in[99:0], 7'h49};
  ZLL_Main_dev8  instR273 (zll_main_dev8_inR73[106:7], zll_main_dev8_inR73[6:0], zll_main_dev8_outR73);
  assign zll_main_dev8_inR74 = {main_dev_in[99:0], 7'h4a};
  ZLL_Main_dev8  instR274 (zll_main_dev8_inR74[106:7], zll_main_dev8_inR74[6:0], zll_main_dev8_outR74);
  assign zll_main_dev8_inR75 = {main_dev_in[99:0], 7'h4b};
  ZLL_Main_dev8  instR275 (zll_main_dev8_inR75[106:7], zll_main_dev8_inR75[6:0], zll_main_dev8_outR75);
  assign zll_main_dev8_inR76 = {main_dev_in[99:0], 7'h4c};
  ZLL_Main_dev8  instR276 (zll_main_dev8_inR76[106:7], zll_main_dev8_inR76[6:0], zll_main_dev8_outR76);
  assign zll_main_dev8_inR77 = {main_dev_in[99:0], 7'h4d};
  ZLL_Main_dev8  instR277 (zll_main_dev8_inR77[106:7], zll_main_dev8_inR77[6:0], zll_main_dev8_outR77);
  assign zll_main_dev8_inR78 = {main_dev_in[99:0], 7'h4e};
  ZLL_Main_dev8  instR278 (zll_main_dev8_inR78[106:7], zll_main_dev8_inR78[6:0], zll_main_dev8_outR78);
  assign zll_main_dev8_inR79 = {main_dev_in[99:0], 7'h4f};
  ZLL_Main_dev8  instR279 (zll_main_dev8_inR79[106:7], zll_main_dev8_inR79[6:0], zll_main_dev8_outR79);
  assign zll_main_dev8_inR80 = {main_dev_in[99:0], 7'h50};
  ZLL_Main_dev8  instR280 (zll_main_dev8_inR80[106:7], zll_main_dev8_inR80[6:0], zll_main_dev8_outR80);
  assign zll_main_dev8_inR81 = {main_dev_in[99:0], 7'h51};
  ZLL_Main_dev8  instR281 (zll_main_dev8_inR81[106:7], zll_main_dev8_inR81[6:0], zll_main_dev8_outR81);
  assign zll_main_dev8_inR82 = {main_dev_in[99:0], 7'h52};
  ZLL_Main_dev8  instR282 (zll_main_dev8_inR82[106:7], zll_main_dev8_inR82[6:0], zll_main_dev8_outR82);
  assign zll_main_dev8_inR83 = {main_dev_in[99:0], 7'h53};
  ZLL_Main_dev8  instR283 (zll_main_dev8_inR83[106:7], zll_main_dev8_inR83[6:0], zll_main_dev8_outR83);
  assign zll_main_dev8_inR84 = {main_dev_in[99:0], 7'h54};
  ZLL_Main_dev8  instR284 (zll_main_dev8_inR84[106:7], zll_main_dev8_inR84[6:0], zll_main_dev8_outR84);
  assign zll_main_dev8_inR85 = {main_dev_in[99:0], 7'h55};
  ZLL_Main_dev8  instR285 (zll_main_dev8_inR85[106:7], zll_main_dev8_inR85[6:0], zll_main_dev8_outR85);
  assign zll_main_dev8_inR86 = {main_dev_in[99:0], 7'h56};
  ZLL_Main_dev8  instR286 (zll_main_dev8_inR86[106:7], zll_main_dev8_inR86[6:0], zll_main_dev8_outR86);
  assign zll_main_dev8_inR87 = {main_dev_in[99:0], 7'h57};
  ZLL_Main_dev8  instR287 (zll_main_dev8_inR87[106:7], zll_main_dev8_inR87[6:0], zll_main_dev8_outR87);
  assign zll_main_dev8_inR88 = {main_dev_in[99:0], 7'h58};
  ZLL_Main_dev8  instR288 (zll_main_dev8_inR88[106:7], zll_main_dev8_inR88[6:0], zll_main_dev8_outR88);
  assign zll_main_dev8_inR89 = {main_dev_in[99:0], 7'h59};
  ZLL_Main_dev8  instR289 (zll_main_dev8_inR89[106:7], zll_main_dev8_inR89[6:0], zll_main_dev8_outR89);
  assign zll_main_dev8_inR90 = {main_dev_in[99:0], 7'h5a};
  ZLL_Main_dev8  instR290 (zll_main_dev8_inR90[106:7], zll_main_dev8_inR90[6:0], zll_main_dev8_outR90);
  assign zll_main_dev8_inR91 = {main_dev_in[99:0], 7'h5b};
  ZLL_Main_dev8  instR291 (zll_main_dev8_inR91[106:7], zll_main_dev8_inR91[6:0], zll_main_dev8_outR91);
  assign zll_main_dev8_inR92 = {main_dev_in[99:0], 7'h5c};
  ZLL_Main_dev8  instR292 (zll_main_dev8_inR92[106:7], zll_main_dev8_inR92[6:0], zll_main_dev8_outR92);
  assign zll_main_dev8_inR93 = {main_dev_in[99:0], 7'h5d};
  ZLL_Main_dev8  instR293 (zll_main_dev8_inR93[106:7], zll_main_dev8_inR93[6:0], zll_main_dev8_outR93);
  assign zll_main_dev8_inR94 = {main_dev_in[99:0], 7'h5e};
  ZLL_Main_dev8  instR294 (zll_main_dev8_inR94[106:7], zll_main_dev8_inR94[6:0], zll_main_dev8_outR94);
  assign zll_main_dev8_inR95 = {main_dev_in[99:0], 7'h5f};
  ZLL_Main_dev8  instR295 (zll_main_dev8_inR95[106:7], zll_main_dev8_inR95[6:0], zll_main_dev8_outR95);
  assign zll_main_dev8_inR96 = {main_dev_in[99:0], 7'h60};
  ZLL_Main_dev8  instR296 (zll_main_dev8_inR96[106:7], zll_main_dev8_inR96[6:0], zll_main_dev8_outR96);
  assign zll_main_dev8_inR97 = {main_dev_in[99:0], 7'h61};
  ZLL_Main_dev8  instR297 (zll_main_dev8_inR97[106:7], zll_main_dev8_inR97[6:0], zll_main_dev8_outR97);
  assign zll_main_dev8_inR98 = {main_dev_in[99:0], 7'h62};
  ZLL_Main_dev8  instR298 (zll_main_dev8_inR98[106:7], zll_main_dev8_inR98[6:0], zll_main_dev8_outR98);
  assign zll_main_dev8_inR99 = {main_dev_in[99:0], 7'h63};
  ZLL_Main_dev8  instR299 (zll_main_dev8_inR99[106:7], zll_main_dev8_inR99[6:0], zll_main_dev8_outR99);
  assign zll_main_dev11_in = {main_dev_in[99:0], 7'h00};
  ZLL_Main_dev11  instR300 (zll_main_dev11_in[106:7], zll_main_dev11_in[6:0], zll_main_dev11_out);
  assign zll_main_dev11_inR1 = {main_dev_in[99:0], 7'h01};
  ZLL_Main_dev11  instR301 (zll_main_dev11_inR1[106:7], zll_main_dev11_inR1[6:0], zll_main_dev11_outR1);
  assign zll_main_dev11_inR2 = {main_dev_in[99:0], 7'h02};
  ZLL_Main_dev11  instR302 (zll_main_dev11_inR2[106:7], zll_main_dev11_inR2[6:0], zll_main_dev11_outR2);
  assign zll_main_dev11_inR3 = {main_dev_in[99:0], 7'h03};
  ZLL_Main_dev11  instR303 (zll_main_dev11_inR3[106:7], zll_main_dev11_inR3[6:0], zll_main_dev11_outR3);
  assign zll_main_dev11_inR4 = {main_dev_in[99:0], 7'h04};
  ZLL_Main_dev11  instR304 (zll_main_dev11_inR4[106:7], zll_main_dev11_inR4[6:0], zll_main_dev11_outR4);
  assign zll_main_dev11_inR5 = {main_dev_in[99:0], 7'h05};
  ZLL_Main_dev11  instR305 (zll_main_dev11_inR5[106:7], zll_main_dev11_inR5[6:0], zll_main_dev11_outR5);
  assign zll_main_dev11_inR6 = {main_dev_in[99:0], 7'h06};
  ZLL_Main_dev11  instR306 (zll_main_dev11_inR6[106:7], zll_main_dev11_inR6[6:0], zll_main_dev11_outR6);
  assign zll_main_dev11_inR7 = {main_dev_in[99:0], 7'h07};
  ZLL_Main_dev11  instR307 (zll_main_dev11_inR7[106:7], zll_main_dev11_inR7[6:0], zll_main_dev11_outR7);
  assign zll_main_dev11_inR8 = {main_dev_in[99:0], 7'h08};
  ZLL_Main_dev11  instR308 (zll_main_dev11_inR8[106:7], zll_main_dev11_inR8[6:0], zll_main_dev11_outR8);
  assign zll_main_dev11_inR9 = {main_dev_in[99:0], 7'h09};
  ZLL_Main_dev11  instR309 (zll_main_dev11_inR9[106:7], zll_main_dev11_inR9[6:0], zll_main_dev11_outR9);
  assign zll_main_dev11_inR10 = {main_dev_in[99:0], 7'h0a};
  ZLL_Main_dev11  instR310 (zll_main_dev11_inR10[106:7], zll_main_dev11_inR10[6:0], zll_main_dev11_outR10);
  assign zll_main_dev11_inR11 = {main_dev_in[99:0], 7'h0b};
  ZLL_Main_dev11  instR311 (zll_main_dev11_inR11[106:7], zll_main_dev11_inR11[6:0], zll_main_dev11_outR11);
  assign zll_main_dev11_inR12 = {main_dev_in[99:0], 7'h0c};
  ZLL_Main_dev11  instR312 (zll_main_dev11_inR12[106:7], zll_main_dev11_inR12[6:0], zll_main_dev11_outR12);
  assign zll_main_dev11_inR13 = {main_dev_in[99:0], 7'h0d};
  ZLL_Main_dev11  instR313 (zll_main_dev11_inR13[106:7], zll_main_dev11_inR13[6:0], zll_main_dev11_outR13);
  assign zll_main_dev11_inR14 = {main_dev_in[99:0], 7'h0e};
  ZLL_Main_dev11  instR314 (zll_main_dev11_inR14[106:7], zll_main_dev11_inR14[6:0], zll_main_dev11_outR14);
  assign zll_main_dev11_inR15 = {main_dev_in[99:0], 7'h0f};
  ZLL_Main_dev11  instR315 (zll_main_dev11_inR15[106:7], zll_main_dev11_inR15[6:0], zll_main_dev11_outR15);
  assign zll_main_dev11_inR16 = {main_dev_in[99:0], 7'h10};
  ZLL_Main_dev11  instR316 (zll_main_dev11_inR16[106:7], zll_main_dev11_inR16[6:0], zll_main_dev11_outR16);
  assign zll_main_dev11_inR17 = {main_dev_in[99:0], 7'h11};
  ZLL_Main_dev11  instR317 (zll_main_dev11_inR17[106:7], zll_main_dev11_inR17[6:0], zll_main_dev11_outR17);
  assign zll_main_dev11_inR18 = {main_dev_in[99:0], 7'h12};
  ZLL_Main_dev11  instR318 (zll_main_dev11_inR18[106:7], zll_main_dev11_inR18[6:0], zll_main_dev11_outR18);
  assign zll_main_dev11_inR19 = {main_dev_in[99:0], 7'h13};
  ZLL_Main_dev11  instR319 (zll_main_dev11_inR19[106:7], zll_main_dev11_inR19[6:0], zll_main_dev11_outR19);
  assign zll_main_dev11_inR20 = {main_dev_in[99:0], 7'h14};
  ZLL_Main_dev11  instR320 (zll_main_dev11_inR20[106:7], zll_main_dev11_inR20[6:0], zll_main_dev11_outR20);
  assign zll_main_dev11_inR21 = {main_dev_in[99:0], 7'h15};
  ZLL_Main_dev11  instR321 (zll_main_dev11_inR21[106:7], zll_main_dev11_inR21[6:0], zll_main_dev11_outR21);
  assign zll_main_dev11_inR22 = {main_dev_in[99:0], 7'h16};
  ZLL_Main_dev11  instR322 (zll_main_dev11_inR22[106:7], zll_main_dev11_inR22[6:0], zll_main_dev11_outR22);
  assign zll_main_dev11_inR23 = {main_dev_in[99:0], 7'h17};
  ZLL_Main_dev11  instR323 (zll_main_dev11_inR23[106:7], zll_main_dev11_inR23[6:0], zll_main_dev11_outR23);
  assign zll_main_dev11_inR24 = {main_dev_in[99:0], 7'h18};
  ZLL_Main_dev11  instR324 (zll_main_dev11_inR24[106:7], zll_main_dev11_inR24[6:0], zll_main_dev11_outR24);
  assign zll_main_dev11_inR25 = {main_dev_in[99:0], 7'h19};
  ZLL_Main_dev11  instR325 (zll_main_dev11_inR25[106:7], zll_main_dev11_inR25[6:0], zll_main_dev11_outR25);
  assign zll_main_dev11_inR26 = {main_dev_in[99:0], 7'h1a};
  ZLL_Main_dev11  instR326 (zll_main_dev11_inR26[106:7], zll_main_dev11_inR26[6:0], zll_main_dev11_outR26);
  assign zll_main_dev11_inR27 = {main_dev_in[99:0], 7'h1b};
  ZLL_Main_dev11  instR327 (zll_main_dev11_inR27[106:7], zll_main_dev11_inR27[6:0], zll_main_dev11_outR27);
  assign zll_main_dev11_inR28 = {main_dev_in[99:0], 7'h1c};
  ZLL_Main_dev11  instR328 (zll_main_dev11_inR28[106:7], zll_main_dev11_inR28[6:0], zll_main_dev11_outR28);
  assign zll_main_dev11_inR29 = {main_dev_in[99:0], 7'h1d};
  ZLL_Main_dev11  instR329 (zll_main_dev11_inR29[106:7], zll_main_dev11_inR29[6:0], zll_main_dev11_outR29);
  assign zll_main_dev11_inR30 = {main_dev_in[99:0], 7'h1e};
  ZLL_Main_dev11  instR330 (zll_main_dev11_inR30[106:7], zll_main_dev11_inR30[6:0], zll_main_dev11_outR30);
  assign zll_main_dev11_inR31 = {main_dev_in[99:0], 7'h1f};
  ZLL_Main_dev11  instR331 (zll_main_dev11_inR31[106:7], zll_main_dev11_inR31[6:0], zll_main_dev11_outR31);
  assign zll_main_dev11_inR32 = {main_dev_in[99:0], 7'h20};
  ZLL_Main_dev11  instR332 (zll_main_dev11_inR32[106:7], zll_main_dev11_inR32[6:0], zll_main_dev11_outR32);
  assign zll_main_dev11_inR33 = {main_dev_in[99:0], 7'h21};
  ZLL_Main_dev11  instR333 (zll_main_dev11_inR33[106:7], zll_main_dev11_inR33[6:0], zll_main_dev11_outR33);
  assign zll_main_dev11_inR34 = {main_dev_in[99:0], 7'h22};
  ZLL_Main_dev11  instR334 (zll_main_dev11_inR34[106:7], zll_main_dev11_inR34[6:0], zll_main_dev11_outR34);
  assign zll_main_dev11_inR35 = {main_dev_in[99:0], 7'h23};
  ZLL_Main_dev11  instR335 (zll_main_dev11_inR35[106:7], zll_main_dev11_inR35[6:0], zll_main_dev11_outR35);
  assign zll_main_dev11_inR36 = {main_dev_in[99:0], 7'h24};
  ZLL_Main_dev11  instR336 (zll_main_dev11_inR36[106:7], zll_main_dev11_inR36[6:0], zll_main_dev11_outR36);
  assign zll_main_dev11_inR37 = {main_dev_in[99:0], 7'h25};
  ZLL_Main_dev11  instR337 (zll_main_dev11_inR37[106:7], zll_main_dev11_inR37[6:0], zll_main_dev11_outR37);
  assign zll_main_dev11_inR38 = {main_dev_in[99:0], 7'h26};
  ZLL_Main_dev11  instR338 (zll_main_dev11_inR38[106:7], zll_main_dev11_inR38[6:0], zll_main_dev11_outR38);
  assign zll_main_dev11_inR39 = {main_dev_in[99:0], 7'h27};
  ZLL_Main_dev11  instR339 (zll_main_dev11_inR39[106:7], zll_main_dev11_inR39[6:0], zll_main_dev11_outR39);
  assign zll_main_dev11_inR40 = {main_dev_in[99:0], 7'h28};
  ZLL_Main_dev11  instR340 (zll_main_dev11_inR40[106:7], zll_main_dev11_inR40[6:0], zll_main_dev11_outR40);
  assign zll_main_dev11_inR41 = {main_dev_in[99:0], 7'h29};
  ZLL_Main_dev11  instR341 (zll_main_dev11_inR41[106:7], zll_main_dev11_inR41[6:0], zll_main_dev11_outR41);
  assign zll_main_dev11_inR42 = {main_dev_in[99:0], 7'h2a};
  ZLL_Main_dev11  instR342 (zll_main_dev11_inR42[106:7], zll_main_dev11_inR42[6:0], zll_main_dev11_outR42);
  assign zll_main_dev11_inR43 = {main_dev_in[99:0], 7'h2b};
  ZLL_Main_dev11  instR343 (zll_main_dev11_inR43[106:7], zll_main_dev11_inR43[6:0], zll_main_dev11_outR43);
  assign zll_main_dev11_inR44 = {main_dev_in[99:0], 7'h2c};
  ZLL_Main_dev11  instR344 (zll_main_dev11_inR44[106:7], zll_main_dev11_inR44[6:0], zll_main_dev11_outR44);
  assign zll_main_dev11_inR45 = {main_dev_in[99:0], 7'h2d};
  ZLL_Main_dev11  instR345 (zll_main_dev11_inR45[106:7], zll_main_dev11_inR45[6:0], zll_main_dev11_outR45);
  assign zll_main_dev11_inR46 = {main_dev_in[99:0], 7'h2e};
  ZLL_Main_dev11  instR346 (zll_main_dev11_inR46[106:7], zll_main_dev11_inR46[6:0], zll_main_dev11_outR46);
  assign zll_main_dev11_inR47 = {main_dev_in[99:0], 7'h2f};
  ZLL_Main_dev11  instR347 (zll_main_dev11_inR47[106:7], zll_main_dev11_inR47[6:0], zll_main_dev11_outR47);
  assign zll_main_dev11_inR48 = {main_dev_in[99:0], 7'h30};
  ZLL_Main_dev11  instR348 (zll_main_dev11_inR48[106:7], zll_main_dev11_inR48[6:0], zll_main_dev11_outR48);
  assign zll_main_dev11_inR49 = {main_dev_in[99:0], 7'h31};
  ZLL_Main_dev11  instR349 (zll_main_dev11_inR49[106:7], zll_main_dev11_inR49[6:0], zll_main_dev11_outR49);
  assign zll_main_dev11_inR50 = {main_dev_in[99:0], 7'h32};
  ZLL_Main_dev11  instR350 (zll_main_dev11_inR50[106:7], zll_main_dev11_inR50[6:0], zll_main_dev11_outR50);
  assign zll_main_dev11_inR51 = {main_dev_in[99:0], 7'h33};
  ZLL_Main_dev11  instR351 (zll_main_dev11_inR51[106:7], zll_main_dev11_inR51[6:0], zll_main_dev11_outR51);
  assign zll_main_dev11_inR52 = {main_dev_in[99:0], 7'h34};
  ZLL_Main_dev11  instR352 (zll_main_dev11_inR52[106:7], zll_main_dev11_inR52[6:0], zll_main_dev11_outR52);
  assign zll_main_dev11_inR53 = {main_dev_in[99:0], 7'h35};
  ZLL_Main_dev11  instR353 (zll_main_dev11_inR53[106:7], zll_main_dev11_inR53[6:0], zll_main_dev11_outR53);
  assign zll_main_dev11_inR54 = {main_dev_in[99:0], 7'h36};
  ZLL_Main_dev11  instR354 (zll_main_dev11_inR54[106:7], zll_main_dev11_inR54[6:0], zll_main_dev11_outR54);
  assign zll_main_dev11_inR55 = {main_dev_in[99:0], 7'h37};
  ZLL_Main_dev11  instR355 (zll_main_dev11_inR55[106:7], zll_main_dev11_inR55[6:0], zll_main_dev11_outR55);
  assign zll_main_dev11_inR56 = {main_dev_in[99:0], 7'h38};
  ZLL_Main_dev11  instR356 (zll_main_dev11_inR56[106:7], zll_main_dev11_inR56[6:0], zll_main_dev11_outR56);
  assign zll_main_dev11_inR57 = {main_dev_in[99:0], 7'h39};
  ZLL_Main_dev11  instR357 (zll_main_dev11_inR57[106:7], zll_main_dev11_inR57[6:0], zll_main_dev11_outR57);
  assign zll_main_dev11_inR58 = {main_dev_in[99:0], 7'h3a};
  ZLL_Main_dev11  instR358 (zll_main_dev11_inR58[106:7], zll_main_dev11_inR58[6:0], zll_main_dev11_outR58);
  assign zll_main_dev11_inR59 = {main_dev_in[99:0], 7'h3b};
  ZLL_Main_dev11  instR359 (zll_main_dev11_inR59[106:7], zll_main_dev11_inR59[6:0], zll_main_dev11_outR59);
  assign zll_main_dev11_inR60 = {main_dev_in[99:0], 7'h3c};
  ZLL_Main_dev11  instR360 (zll_main_dev11_inR60[106:7], zll_main_dev11_inR60[6:0], zll_main_dev11_outR60);
  assign zll_main_dev11_inR61 = {main_dev_in[99:0], 7'h3d};
  ZLL_Main_dev11  instR361 (zll_main_dev11_inR61[106:7], zll_main_dev11_inR61[6:0], zll_main_dev11_outR61);
  assign zll_main_dev11_inR62 = {main_dev_in[99:0], 7'h3e};
  ZLL_Main_dev11  instR362 (zll_main_dev11_inR62[106:7], zll_main_dev11_inR62[6:0], zll_main_dev11_outR62);
  assign zll_main_dev11_inR63 = {main_dev_in[99:0], 7'h3f};
  ZLL_Main_dev11  instR363 (zll_main_dev11_inR63[106:7], zll_main_dev11_inR63[6:0], zll_main_dev11_outR63);
  assign zll_main_dev11_inR64 = {main_dev_in[99:0], 7'h40};
  ZLL_Main_dev11  instR364 (zll_main_dev11_inR64[106:7], zll_main_dev11_inR64[6:0], zll_main_dev11_outR64);
  assign zll_main_dev11_inR65 = {main_dev_in[99:0], 7'h41};
  ZLL_Main_dev11  instR365 (zll_main_dev11_inR65[106:7], zll_main_dev11_inR65[6:0], zll_main_dev11_outR65);
  assign zll_main_dev11_inR66 = {main_dev_in[99:0], 7'h42};
  ZLL_Main_dev11  instR366 (zll_main_dev11_inR66[106:7], zll_main_dev11_inR66[6:0], zll_main_dev11_outR66);
  assign zll_main_dev11_inR67 = {main_dev_in[99:0], 7'h43};
  ZLL_Main_dev11  instR367 (zll_main_dev11_inR67[106:7], zll_main_dev11_inR67[6:0], zll_main_dev11_outR67);
  assign zll_main_dev11_inR68 = {main_dev_in[99:0], 7'h44};
  ZLL_Main_dev11  instR368 (zll_main_dev11_inR68[106:7], zll_main_dev11_inR68[6:0], zll_main_dev11_outR68);
  assign zll_main_dev11_inR69 = {main_dev_in[99:0], 7'h45};
  ZLL_Main_dev11  instR369 (zll_main_dev11_inR69[106:7], zll_main_dev11_inR69[6:0], zll_main_dev11_outR69);
  assign zll_main_dev11_inR70 = {main_dev_in[99:0], 7'h46};
  ZLL_Main_dev11  instR370 (zll_main_dev11_inR70[106:7], zll_main_dev11_inR70[6:0], zll_main_dev11_outR70);
  assign zll_main_dev11_inR71 = {main_dev_in[99:0], 7'h47};
  ZLL_Main_dev11  instR371 (zll_main_dev11_inR71[106:7], zll_main_dev11_inR71[6:0], zll_main_dev11_outR71);
  assign zll_main_dev11_inR72 = {main_dev_in[99:0], 7'h48};
  ZLL_Main_dev11  instR372 (zll_main_dev11_inR72[106:7], zll_main_dev11_inR72[6:0], zll_main_dev11_outR72);
  assign zll_main_dev11_inR73 = {main_dev_in[99:0], 7'h49};
  ZLL_Main_dev11  instR373 (zll_main_dev11_inR73[106:7], zll_main_dev11_inR73[6:0], zll_main_dev11_outR73);
  assign zll_main_dev11_inR74 = {main_dev_in[99:0], 7'h4a};
  ZLL_Main_dev11  instR374 (zll_main_dev11_inR74[106:7], zll_main_dev11_inR74[6:0], zll_main_dev11_outR74);
  assign zll_main_dev11_inR75 = {main_dev_in[99:0], 7'h4b};
  ZLL_Main_dev11  instR375 (zll_main_dev11_inR75[106:7], zll_main_dev11_inR75[6:0], zll_main_dev11_outR75);
  assign zll_main_dev11_inR76 = {main_dev_in[99:0], 7'h4c};
  ZLL_Main_dev11  instR376 (zll_main_dev11_inR76[106:7], zll_main_dev11_inR76[6:0], zll_main_dev11_outR76);
  assign zll_main_dev11_inR77 = {main_dev_in[99:0], 7'h4d};
  ZLL_Main_dev11  instR377 (zll_main_dev11_inR77[106:7], zll_main_dev11_inR77[6:0], zll_main_dev11_outR77);
  assign zll_main_dev11_inR78 = {main_dev_in[99:0], 7'h4e};
  ZLL_Main_dev11  instR378 (zll_main_dev11_inR78[106:7], zll_main_dev11_inR78[6:0], zll_main_dev11_outR78);
  assign zll_main_dev11_inR79 = {main_dev_in[99:0], 7'h4f};
  ZLL_Main_dev11  instR379 (zll_main_dev11_inR79[106:7], zll_main_dev11_inR79[6:0], zll_main_dev11_outR79);
  assign zll_main_dev11_inR80 = {main_dev_in[99:0], 7'h50};
  ZLL_Main_dev11  instR380 (zll_main_dev11_inR80[106:7], zll_main_dev11_inR80[6:0], zll_main_dev11_outR80);
  assign zll_main_dev11_inR81 = {main_dev_in[99:0], 7'h51};
  ZLL_Main_dev11  instR381 (zll_main_dev11_inR81[106:7], zll_main_dev11_inR81[6:0], zll_main_dev11_outR81);
  assign zll_main_dev11_inR82 = {main_dev_in[99:0], 7'h52};
  ZLL_Main_dev11  instR382 (zll_main_dev11_inR82[106:7], zll_main_dev11_inR82[6:0], zll_main_dev11_outR82);
  assign zll_main_dev11_inR83 = {main_dev_in[99:0], 7'h53};
  ZLL_Main_dev11  instR383 (zll_main_dev11_inR83[106:7], zll_main_dev11_inR83[6:0], zll_main_dev11_outR83);
  assign zll_main_dev11_inR84 = {main_dev_in[99:0], 7'h54};
  ZLL_Main_dev11  instR384 (zll_main_dev11_inR84[106:7], zll_main_dev11_inR84[6:0], zll_main_dev11_outR84);
  assign zll_main_dev11_inR85 = {main_dev_in[99:0], 7'h55};
  ZLL_Main_dev11  instR385 (zll_main_dev11_inR85[106:7], zll_main_dev11_inR85[6:0], zll_main_dev11_outR85);
  assign zll_main_dev11_inR86 = {main_dev_in[99:0], 7'h56};
  ZLL_Main_dev11  instR386 (zll_main_dev11_inR86[106:7], zll_main_dev11_inR86[6:0], zll_main_dev11_outR86);
  assign zll_main_dev11_inR87 = {main_dev_in[99:0], 7'h57};
  ZLL_Main_dev11  instR387 (zll_main_dev11_inR87[106:7], zll_main_dev11_inR87[6:0], zll_main_dev11_outR87);
  assign zll_main_dev11_inR88 = {main_dev_in[99:0], 7'h58};
  ZLL_Main_dev11  instR388 (zll_main_dev11_inR88[106:7], zll_main_dev11_inR88[6:0], zll_main_dev11_outR88);
  assign zll_main_dev11_inR89 = {main_dev_in[99:0], 7'h59};
  ZLL_Main_dev11  instR389 (zll_main_dev11_inR89[106:7], zll_main_dev11_inR89[6:0], zll_main_dev11_outR89);
  assign zll_main_dev11_inR90 = {main_dev_in[99:0], 7'h5a};
  ZLL_Main_dev11  instR390 (zll_main_dev11_inR90[106:7], zll_main_dev11_inR90[6:0], zll_main_dev11_outR90);
  assign zll_main_dev11_inR91 = {main_dev_in[99:0], 7'h5b};
  ZLL_Main_dev11  instR391 (zll_main_dev11_inR91[106:7], zll_main_dev11_inR91[6:0], zll_main_dev11_outR91);
  assign zll_main_dev11_inR92 = {main_dev_in[99:0], 7'h5c};
  ZLL_Main_dev11  instR392 (zll_main_dev11_inR92[106:7], zll_main_dev11_inR92[6:0], zll_main_dev11_outR92);
  assign zll_main_dev11_inR93 = {main_dev_in[99:0], 7'h5d};
  ZLL_Main_dev11  instR393 (zll_main_dev11_inR93[106:7], zll_main_dev11_inR93[6:0], zll_main_dev11_outR93);
  assign zll_main_dev11_inR94 = {main_dev_in[99:0], 7'h5e};
  ZLL_Main_dev11  instR394 (zll_main_dev11_inR94[106:7], zll_main_dev11_inR94[6:0], zll_main_dev11_outR94);
  assign zll_main_dev11_inR95 = {main_dev_in[99:0], 7'h5f};
  ZLL_Main_dev11  instR395 (zll_main_dev11_inR95[106:7], zll_main_dev11_inR95[6:0], zll_main_dev11_outR95);
  assign zll_main_dev11_inR96 = {main_dev_in[99:0], 7'h60};
  ZLL_Main_dev11  instR396 (zll_main_dev11_inR96[106:7], zll_main_dev11_inR96[6:0], zll_main_dev11_outR96);
  assign zll_main_dev11_inR97 = {main_dev_in[99:0], 7'h61};
  ZLL_Main_dev11  instR397 (zll_main_dev11_inR97[106:7], zll_main_dev11_inR97[6:0], zll_main_dev11_outR97);
  assign zll_main_dev11_inR98 = {main_dev_in[99:0], 7'h62};
  ZLL_Main_dev11  instR398 (zll_main_dev11_inR98[106:7], zll_main_dev11_inR98[6:0], zll_main_dev11_outR98);
  assign zll_main_dev11_inR99 = {main_dev_in[99:0], 7'h63};
  ZLL_Main_dev11  instR399 (zll_main_dev11_inR99[106:7], zll_main_dev11_inR99[6:0], zll_main_dev11_outR99);
  assign {__continue, __out0, __out1, __out2, __out3, __resumption_tag_next} = {zll_main_dev2_out, zll_main_dev2_outR1, zll_main_dev2_outR2, zll_main_dev2_outR3, zll_main_dev2_outR4, zll_main_dev2_outR5, zll_main_dev2_outR6, zll_main_dev2_outR7, zll_main_dev2_outR8, zll_main_dev2_outR9, zll_main_dev2_outR10, zll_main_dev2_outR11, zll_main_dev2_outR12, zll_main_dev2_outR13, zll_main_dev2_outR14, zll_main_dev2_outR15, zll_main_dev2_outR16, zll_main_dev2_outR17, zll_main_dev2_outR18, zll_main_dev2_outR19, zll_main_dev2_outR20, zll_main_dev2_outR21, zll_main_dev2_outR22, zll_main_dev2_outR23, zll_main_dev2_outR24, zll_main_dev2_outR25, zll_main_dev2_outR26, zll_main_dev2_outR27, zll_main_dev2_outR28, zll_main_dev2_outR29, zll_main_dev2_outR30, zll_main_dev2_outR31, zll_main_dev2_outR32, zll_main_dev2_outR33, zll_main_dev2_outR34, zll_main_dev2_outR35, zll_main_dev2_outR36, zll_main_dev2_outR37, zll_main_dev2_outR38, zll_main_dev2_outR39, zll_main_dev2_outR40, zll_main_dev2_outR41, zll_main_dev2_outR42, zll_main_dev2_outR43, zll_main_dev2_outR44, zll_main_dev2_outR45, zll_main_dev2_outR46, zll_main_dev2_outR47, zll_main_dev2_outR48, zll_main_dev2_outR49, zll_main_dev2_outR50, zll_main_dev2_outR51, zll_main_dev2_outR52, zll_main_dev2_outR53, zll_main_dev2_outR54, zll_main_dev2_outR55, zll_main_dev2_outR56, zll_main_dev2_outR57, zll_main_dev2_outR58, zll_main_dev2_outR59, zll_main_dev2_outR60, zll_main_dev2_outR61, zll_main_dev2_outR62, zll_main_dev2_outR63, zll_main_dev2_outR64, zll_main_dev2_outR65, zll_main_dev2_outR66, zll_main_dev2_outR67, zll_main_dev2_outR68, zll_main_dev2_outR69, zll_main_dev2_outR70, zll_main_dev2_outR71, zll_main_dev2_outR72, zll_main_dev2_outR73, zll_main_dev2_outR74, zll_main_dev2_outR75, zll_main_dev2_outR76, zll_main_dev2_outR77, zll_main_dev2_outR78, zll_main_dev2_outR79, zll_main_dev2_outR80, zll_main_dev2_outR81, zll_main_dev2_outR82, zll_main_dev2_outR83, zll_main_dev2_outR84, zll_main_dev2_outR85, zll_main_dev2_outR86, zll_main_dev2_outR87, zll_main_dev2_outR88, zll_main_dev2_outR89, zll_main_dev2_outR90, zll_main_dev2_outR91, zll_main_dev2_outR92, zll_main_dev2_outR93, zll_main_dev2_outR94, zll_main_dev2_outR95, zll_main_dev2_outR96, zll_main_dev2_outR97, zll_main_dev2_outR98, zll_main_dev2_outR99, zll_main_dev5_out, zll_main_dev5_outR1, zll_main_dev5_outR2, zll_main_dev5_outR3, zll_main_dev5_outR4, zll_main_dev5_outR5, zll_main_dev5_outR6, zll_main_dev5_outR7, zll_main_dev5_outR8, zll_main_dev5_outR9, zll_main_dev5_outR10, zll_main_dev5_outR11, zll_main_dev5_outR12, zll_main_dev5_outR13, zll_main_dev5_outR14, zll_main_dev5_outR15, zll_main_dev5_outR16, zll_main_dev5_outR17, zll_main_dev5_outR18, zll_main_dev5_outR19, zll_main_dev5_outR20, zll_main_dev5_outR21, zll_main_dev5_outR22, zll_main_dev5_outR23, zll_main_dev5_outR24, zll_main_dev5_outR25, zll_main_dev5_outR26, zll_main_dev5_outR27, zll_main_dev5_outR28, zll_main_dev5_outR29, zll_main_dev5_outR30, zll_main_dev5_outR31, zll_main_dev5_outR32, zll_main_dev5_outR33, zll_main_dev5_outR34, zll_main_dev5_outR35, zll_main_dev5_outR36, zll_main_dev5_outR37, zll_main_dev5_outR38, zll_main_dev5_outR39, zll_main_dev5_outR40, zll_main_dev5_outR41, zll_main_dev5_outR42, zll_main_dev5_outR43, zll_main_dev5_outR44, zll_main_dev5_outR45, zll_main_dev5_outR46, zll_main_dev5_outR47, zll_main_dev5_outR48, zll_main_dev5_outR49, zll_main_dev5_outR50, zll_main_dev5_outR51, zll_main_dev5_outR52, zll_main_dev5_outR53, zll_main_dev5_outR54, zll_main_dev5_outR55, zll_main_dev5_outR56, zll_main_dev5_outR57, zll_main_dev5_outR58, zll_main_dev5_outR59, zll_main_dev5_outR60, zll_main_dev5_outR61, zll_main_dev5_outR62, zll_main_dev5_outR63, zll_main_dev5_outR64, zll_main_dev5_outR65, zll_main_dev5_outR66, zll_main_dev5_outR67, zll_main_dev5_outR68, zll_main_dev5_outR69, zll_main_dev5_outR70, zll_main_dev5_outR71, zll_main_dev5_outR72, zll_main_dev5_outR73, zll_main_dev5_outR74, zll_main_dev5_outR75, zll_main_dev5_outR76, zll_main_dev5_outR77, zll_main_dev5_outR78, zll_main_dev5_outR79, zll_main_dev5_outR80, zll_main_dev5_outR81, zll_main_dev5_outR82, zll_main_dev5_outR83, zll_main_dev5_outR84, zll_main_dev5_outR85, zll_main_dev5_outR86, zll_main_dev5_outR87, zll_main_dev5_outR88, zll_main_dev5_outR89, zll_main_dev5_outR90, zll_main_dev5_outR91, zll_main_dev5_outR92, zll_main_dev5_outR93, zll_main_dev5_outR94, zll_main_dev5_outR95, zll_main_dev5_outR96, zll_main_dev5_outR97, zll_main_dev5_outR98, zll_main_dev5_outR99, zll_main_dev8_out, zll_main_dev8_outR1, zll_main_dev8_outR2, zll_main_dev8_outR3, zll_main_dev8_outR4, zll_main_dev8_outR5, zll_main_dev8_outR6, zll_main_dev8_outR7, zll_main_dev8_outR8, zll_main_dev8_outR9, zll_main_dev8_outR10, zll_main_dev8_outR11, zll_main_dev8_outR12, zll_main_dev8_outR13, zll_main_dev8_outR14, zll_main_dev8_outR15, zll_main_dev8_outR16, zll_main_dev8_outR17, zll_main_dev8_outR18, zll_main_dev8_outR19, zll_main_dev8_outR20, zll_main_dev8_outR21, zll_main_dev8_outR22, zll_main_dev8_outR23, zll_main_dev8_outR24, zll_main_dev8_outR25, zll_main_dev8_outR26, zll_main_dev8_outR27, zll_main_dev8_outR28, zll_main_dev8_outR29, zll_main_dev8_outR30, zll_main_dev8_outR31, zll_main_dev8_outR32, zll_main_dev8_outR33, zll_main_dev8_outR34, zll_main_dev8_outR35, zll_main_dev8_outR36, zll_main_dev8_outR37, zll_main_dev8_outR38, zll_main_dev8_outR39, zll_main_dev8_outR40, zll_main_dev8_outR41, zll_main_dev8_outR42, zll_main_dev8_outR43, zll_main_dev8_outR44, zll_main_dev8_outR45, zll_main_dev8_outR46, zll_main_dev8_outR47, zll_main_dev8_outR48, zll_main_dev8_outR49, zll_main_dev8_outR50, zll_main_dev8_outR51, zll_main_dev8_outR52, zll_main_dev8_outR53, zll_main_dev8_outR54, zll_main_dev8_outR55, zll_main_dev8_outR56, zll_main_dev8_outR57, zll_main_dev8_outR58, zll_main_dev8_outR59, zll_main_dev8_outR60, zll_main_dev8_outR61, zll_main_dev8_outR62, zll_main_dev8_outR63, zll_main_dev8_outR64, zll_main_dev8_outR65, zll_main_dev8_outR66, zll_main_dev8_outR67, zll_main_dev8_outR68, zll_main_dev8_outR69, zll_main_dev8_outR70, zll_main_dev8_outR71, zll_main_dev8_outR72, zll_main_dev8_outR73, zll_main_dev8_outR74, zll_main_dev8_outR75, zll_main_dev8_outR76, zll_main_dev8_outR77, zll_main_dev8_outR78, zll_main_dev8_outR79, zll_main_dev8_outR80, zll_main_dev8_outR81, zll_main_dev8_outR82, zll_main_dev8_outR83, zll_main_dev8_outR84, zll_main_dev8_outR85, zll_main_dev8_outR86, zll_main_dev8_outR87, zll_main_dev8_outR88, zll_main_dev8_outR89, zll_main_dev8_outR90, zll_main_dev8_outR91, zll_main_dev8_outR92, zll_main_dev8_outR93, zll_main_dev8_outR94, zll_main_dev8_outR95, zll_main_dev8_outR96, zll_main_dev8_outR97, zll_main_dev8_outR98, zll_main_dev8_outR99, zll_main_dev11_out, zll_main_dev11_outR1, zll_main_dev11_outR2, zll_main_dev11_outR3, zll_main_dev11_outR4, zll_main_dev11_outR5, zll_main_dev11_outR6, zll_main_dev11_outR7, zll_main_dev11_outR8, zll_main_dev11_outR9, zll_main_dev11_outR10, zll_main_dev11_outR11, zll_main_dev11_outR12, zll_main_dev11_outR13, zll_main_dev11_outR14, zll_main_dev11_outR15, zll_main_dev11_outR16, zll_main_dev11_outR17, zll_main_dev11_outR18, zll_main_dev11_outR19, zll_main_dev11_outR20, zll_main_dev11_outR21, zll_main_dev11_outR22, zll_main_dev11_outR23, zll_main_dev11_outR24, zll_main_dev11_outR25, zll_main_dev11_outR26, zll_main_dev11_outR27, zll_main_dev11_outR28, zll_main_dev11_outR29, zll_main_dev11_outR30, zll_main_dev11_outR31, zll_main_dev11_outR32, zll_main_dev11_outR33, zll_main_dev11_outR34, zll_main_dev11_outR35, zll_main_dev11_outR36, zll_main_dev11_outR37, zll_main_dev11_outR38, zll_main_dev11_outR39, zll_main_dev11_outR40, zll_main_dev11_outR41, zll_main_dev11_outR42, zll_main_dev11_outR43, zll_main_dev11_outR44, zll_main_dev11_outR45, zll_main_dev11_outR46, zll_main_dev11_outR47, zll_main_dev11_outR48, zll_main_dev11_outR49, zll_main_dev11_outR50, zll_main_dev11_outR51, zll_main_dev11_outR52, zll_main_dev11_outR53, zll_main_dev11_outR54, zll_main_dev11_outR55, zll_main_dev11_outR56, zll_main_dev11_outR57, zll_main_dev11_outR58, zll_main_dev11_outR59, zll_main_dev11_outR60, zll_main_dev11_outR61, zll_main_dev11_outR62, zll_main_dev11_outR63, zll_main_dev11_outR64, zll_main_dev11_outR65, zll_main_dev11_outR66, zll_main_dev11_outR67, zll_main_dev11_outR68, zll_main_dev11_outR69, zll_main_dev11_outR70, zll_main_dev11_outR71, zll_main_dev11_outR72, zll_main_dev11_outR73, zll_main_dev11_outR74, zll_main_dev11_outR75, zll_main_dev11_outR76, zll_main_dev11_outR77, zll_main_dev11_outR78, zll_main_dev11_outR79, zll_main_dev11_outR80, zll_main_dev11_outR81, zll_main_dev11_outR82, zll_main_dev11_outR83, zll_main_dev11_outR84, zll_main_dev11_outR85, zll_main_dev11_outR86, zll_main_dev11_outR87, zll_main_dev11_outR88, zll_main_dev11_outR89, zll_main_dev11_outR90, zll_main_dev11_outR91, zll_main_dev11_outR92, zll_main_dev11_outR93, zll_main_dev11_outR94, zll_main_dev11_outR95, zll_main_dev11_outR96, zll_main_dev11_outR97, zll_main_dev11_outR98, zll_main_dev11_outR99};
  initial __resumption_tag <= {7'h64{1'h0}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      __resumption_tag <= {7'h64{1'h0}};
    end else begin
      __resumption_tag <= __resumption_tag_next;
    end
  end
endmodule

module ZLL_Main_dev2 (input logic [99:0] arg0,
  input logic [6:0] arg1,
  output logic [0:0] res);
  logic [6:0] resize_in;
  logic [127:0] resize_inR1;
  logic [0:0] msbit_in;
  logic [0:0] rewire_prelude_not_in;
  logic [0:0] rewire_prelude_not_out;
  logic [6:0] resize_inR2;
  logic [127:0] resize_inR3;
  logic [0:0] msbit_inR1;
  logic [0:0] rewire_prelude_not_inR1;
  logic [0:0] rewire_prelude_not_outR1;
  logic [107:0] zll_main_dev1_in;
  logic [99:0] main_x2_in;
  logic [99:0] main_x2_out;
  logic [99:0] resize_inR4;
  logic [6:0] resize_inR5;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR6;
  logic [6:0] resize_inR7;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR8;
  logic [6:0] resize_inR9;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR10;
  logic [107:0] zll_main_dev_in;
  logic [99:0] resize_inR11;
  logic [6:0] resize_inR12;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR13;
  logic [6:0] resize_inR14;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [127:0] resize_inR15;
  assign resize_in = arg1;
  assign resize_inR1 = 128'(resize_in[6:0]);
  assign msbit_in = resize_inR1[0];
  assign rewire_prelude_not_in = msbit_in[0];
  ReWire_Prelude_not  inst (rewire_prelude_not_in[0], rewire_prelude_not_out);
  assign resize_inR2 = arg1;
  assign resize_inR3 = 128'(resize_inR2[6:0]);
  assign msbit_inR1 = resize_inR3[0];
  assign rewire_prelude_not_inR1 = msbit_inR1[0];
  ReWire_Prelude_not  instR1 (rewire_prelude_not_inR1[0], rewire_prelude_not_outR1);
  assign zll_main_dev1_in = {arg0, arg1, rewire_prelude_not_outR1};
  assign main_x2_in = zll_main_dev1_in[107:8];
  Main_x2  instR2 (main_x2_in[99:0], main_x2_out);
  assign resize_inR4 = main_x2_out;
  assign resize_inR5 = zll_main_dev1_in[7:1];
  assign binop_in = {128'(resize_inR5[6:0]), 128'h00000000000000000000000000000001};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h00000000000000000000000000000064};
  assign resize_inR6 = binop_inR1[255:128] % binop_inR1[127:0];
  assign resize_inR7 = resize_inR6[6:0];
  assign binop_inR2 = {128'(resize_inR7[6:0]), 128'h00000000000000000000000000000002};
  assign binop_inR3 = {binop_inR2[255:128] / binop_inR2[127:0], 128'h00000000000000000000000000000064};
  assign resize_inR8 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR9 = resize_inR8[6:0];
  assign binop_inR4 = {128'h00000000000000000000000000000064, 128'(resize_inR9[6:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR7 = {128'(resize_inR4[99:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR10 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign zll_main_dev_in = {arg0, arg1, rewire_prelude_not_out};
  assign resize_inR11 = zll_main_dev_in[107:8];
  assign resize_inR12 = zll_main_dev_in[7:1];
  assign binop_inR8 = {128'(resize_inR12[6:0]), 128'h00000000000000000000000000000002};
  assign binop_inR9 = {binop_inR8[255:128] / binop_inR8[127:0], 128'h00000000000000000000000000000064};
  assign resize_inR13 = binop_inR9[255:128] % binop_inR9[127:0];
  assign resize_inR14 = resize_inR13[6:0];
  assign binop_inR10 = {128'h00000000000000000000000000000064, 128'(resize_inR14[6:0])};
  assign binop_inR11 = {binop_inR10[255:128] - binop_inR10[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR12 = {binop_inR11[255:128] - binop_inR11[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR13 = {128'(resize_inR11[99:0]), binop_inR12[255:128] * binop_inR12[127:0]};
  assign resize_inR15 = binop_inR13[255:128] >> binop_inR13[127:0];
  assign res = (zll_main_dev_in[0] == 1'h1) ? resize_inR15[0] : resize_inR10[0];
endmodule

module ZLL_Main_dev5 (input logic [99:0] arg0,
  input logic [6:0] arg1,
  output logic [0:0] res);
  logic [6:0] resize_in;
  logic [127:0] resize_inR1;
  logic [0:0] msbit_in;
  logic [0:0] rewire_prelude_not_in;
  logic [0:0] rewire_prelude_not_out;
  logic [6:0] resize_inR2;
  logic [127:0] resize_inR3;
  logic [0:0] msbit_inR1;
  logic [0:0] rewire_prelude_not_inR1;
  logic [0:0] rewire_prelude_not_outR1;
  logic [107:0] zll_main_dev4_in;
  logic [99:0] main_x2_in;
  logic [99:0] main_x2_out;
  logic [99:0] resize_inR4;
  logic [6:0] resize_inR5;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR6;
  logic [6:0] resize_inR7;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR8;
  logic [6:0] resize_inR9;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR10;
  logic [6:0] resize_inR11;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR12;
  logic [107:0] zll_main_dev3_in;
  logic [99:0] resize_inR13;
  logic [6:0] resize_inR14;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR15;
  logic [6:0] resize_inR16;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [127:0] resize_inR17;
  logic [6:0] resize_inR18;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [255:0] binop_inR16;
  logic [255:0] binop_inR17;
  logic [127:0] resize_inR19;
  assign resize_in = arg1;
  assign resize_inR1 = 128'(resize_in[6:0]);
  assign msbit_in = resize_inR1[0];
  assign rewire_prelude_not_in = msbit_in[0];
  ReWire_Prelude_not  inst (rewire_prelude_not_in[0], rewire_prelude_not_out);
  assign resize_inR2 = arg1;
  assign resize_inR3 = 128'(resize_inR2[6:0]);
  assign msbit_inR1 = resize_inR3[0];
  assign rewire_prelude_not_inR1 = msbit_inR1[0];
  ReWire_Prelude_not  instR1 (rewire_prelude_not_inR1[0], rewire_prelude_not_outR1);
  assign zll_main_dev4_in = {arg0, arg1, rewire_prelude_not_outR1};
  assign main_x2_in = zll_main_dev4_in[107:8];
  Main_x2  instR2 (main_x2_in[99:0], main_x2_out);
  assign resize_inR4 = main_x2_out;
  assign resize_inR5 = zll_main_dev4_in[7:1];
  assign binop_in = {128'(resize_inR5[6:0]), 128'h00000000000000000000000000000001};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h00000000000000000000000000000064};
  assign resize_inR6 = binop_inR1[255:128] % binop_inR1[127:0];
  assign resize_inR7 = resize_inR6[6:0];
  assign binop_inR2 = {128'h00000000000000000000000000000031, 128'(resize_inR7[6:0])};
  assign binop_inR3 = {binop_inR2[255:128] + binop_inR2[127:0], 128'h00000000000000000000000000000064};
  assign resize_inR8 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR9 = resize_inR8[6:0];
  assign binop_inR4 = {128'(resize_inR9[6:0]), 128'h00000000000000000000000000000002};
  assign binop_inR5 = {binop_inR4[255:128] / binop_inR4[127:0], 128'h00000000000000000000000000000064};
  assign resize_inR10 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR11 = resize_inR10[6:0];
  assign binop_inR6 = {128'h00000000000000000000000000000064, 128'(resize_inR11[6:0])};
  assign binop_inR7 = {binop_inR6[255:128] - binop_inR6[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR8 = {binop_inR7[255:128] - binop_inR7[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR9 = {128'(resize_inR4[99:0]), binop_inR8[255:128] * binop_inR8[127:0]};
  assign resize_inR12 = binop_inR9[255:128] >> binop_inR9[127:0];
  assign zll_main_dev3_in = {arg0, arg1, rewire_prelude_not_out};
  assign resize_inR13 = zll_main_dev3_in[107:8];
  assign resize_inR14 = zll_main_dev3_in[7:1];
  assign binop_inR10 = {128'h00000000000000000000000000000031, 128'(resize_inR14[6:0])};
  assign binop_inR11 = {binop_inR10[255:128] + binop_inR10[127:0], 128'h00000000000000000000000000000064};
  assign resize_inR15 = binop_inR11[255:128] % binop_inR11[127:0];
  assign resize_inR16 = resize_inR15[6:0];
  assign binop_inR12 = {128'(resize_inR16[6:0]), 128'h00000000000000000000000000000002};
  assign binop_inR13 = {binop_inR12[255:128] / binop_inR12[127:0], 128'h00000000000000000000000000000064};
  assign resize_inR17 = binop_inR13[255:128] % binop_inR13[127:0];
  assign resize_inR18 = resize_inR17[6:0];
  assign binop_inR14 = {128'h00000000000000000000000000000064, 128'(resize_inR18[6:0])};
  assign binop_inR15 = {binop_inR14[255:128] - binop_inR14[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR16 = {binop_inR15[255:128] - binop_inR15[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR17 = {128'(resize_inR13[99:0]), binop_inR16[255:128] * binop_inR16[127:0]};
  assign resize_inR19 = binop_inR17[255:128] >> binop_inR17[127:0];
  assign res = (zll_main_dev3_in[0] == 1'h1) ? resize_inR19[0] : resize_inR12[0];
endmodule

module ZLL_Main_dev8 (input logic [99:0] arg0,
  input logic [6:0] arg1,
  output logic [0:0] res);
  logic [6:0] resize_in;
  logic [255:0] binop_in;
  logic [6:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [107:0] zll_main_dev7_in;
  logic [99:0] main_x2_in;
  logic [99:0] main_x2_out;
  logic [99:0] resize_inR2;
  logic [6:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [6:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [6:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR8;
  logic [107:0] zll_main_dev6_in;
  logic [99:0] resize_inR9;
  logic [6:0] resize_inR10;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR11;
  logic [6:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR13;
  assign resize_in = arg1;
  assign binop_in = {128'(resize_in[6:0]), 128'h00000000000000000000000000000031};
  assign resize_inR1 = arg1;
  assign binop_inR1 = {128'(resize_inR1[6:0]), 128'h00000000000000000000000000000031};
  assign zll_main_dev7_in = {arg0, arg1, binop_inR1[255:128] < binop_inR1[127:0]};
  assign main_x2_in = zll_main_dev7_in[107:8];
  Main_x2  inst (main_x2_in[99:0], main_x2_out);
  assign resize_inR2 = main_x2_out;
  assign resize_inR3 = zll_main_dev7_in[7:1];
  assign binop_inR2 = {128'(resize_inR3[6:0]), 128'h00000000000000000000000000000031};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h00000000000000000000000000000064};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[6:0];
  assign binop_inR4 = {128'(resize_inR5[6:0]), 128'h00000000000000000000000000000002};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h00000000000000000000000000000064};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[6:0];
  assign binop_inR6 = {128'h00000000000000000000000000000064, 128'(resize_inR7[6:0])};
  assign binop_inR7 = {binop_inR6[255:128] - binop_inR6[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR8 = {binop_inR7[255:128] - binop_inR7[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR9 = {128'(resize_inR2[99:0]), binop_inR8[255:128] * binop_inR8[127:0]};
  assign resize_inR8 = binop_inR9[255:128] >> binop_inR9[127:0];
  assign zll_main_dev6_in = {arg0, arg1, binop_in[255:128] < binop_in[127:0]};
  assign resize_inR9 = zll_main_dev6_in[107:8];
  assign resize_inR10 = zll_main_dev6_in[7:1];
  assign binop_inR10 = {128'(resize_inR10[6:0]), 128'h00000000000000000000000000000002};
  assign binop_inR11 = {binop_inR10[255:128] * binop_inR10[127:0], 128'h00000000000000000000000000000064};
  assign resize_inR11 = binop_inR11[255:128] % binop_inR11[127:0];
  assign resize_inR12 = resize_inR11[6:0];
  assign binop_inR12 = {128'h00000000000000000000000000000064, 128'(resize_inR12[6:0])};
  assign binop_inR13 = {binop_inR12[255:128] - binop_inR12[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR14 = {binop_inR13[255:128] - binop_inR13[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR15 = {128'(resize_inR9[99:0]), binop_inR14[255:128] * binop_inR14[127:0]};
  assign resize_inR13 = binop_inR15[255:128] >> binop_inR15[127:0];
  assign res = (zll_main_dev6_in[0] == 1'h1) ? resize_inR13[0] : resize_inR8[0];
endmodule

module ZLL_Main_dev11 (input logic [99:0] arg0,
  input logic [6:0] arg1,
  output logic [0:0] res);
  logic [6:0] resize_in;
  logic [255:0] binop_in;
  logic [6:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [107:0] zll_main_dev10_in;
  logic [99:0] main_x2_in;
  logic [99:0] main_x2_out;
  logic [99:0] resize_inR2;
  logic [6:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [6:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [6:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR8;
  logic [6:0] resize_inR9;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR10;
  logic [107:0] zll_main_dev9_in;
  logic [99:0] resize_inR11;
  logic [6:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [127:0] resize_inR13;
  logic [6:0] resize_inR14;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR15;
  logic [6:0] resize_inR16;
  logic [255:0] binop_inR16;
  logic [255:0] binop_inR17;
  logic [255:0] binop_inR18;
  logic [255:0] binop_inR19;
  logic [127:0] resize_inR17;
  assign resize_in = arg1;
  assign binop_in = {128'(resize_in[6:0]), 128'h00000000000000000000000000000031};
  assign resize_inR1 = arg1;
  assign binop_inR1 = {128'(resize_inR1[6:0]), 128'h00000000000000000000000000000031};
  assign zll_main_dev10_in = {arg0, arg1, binop_inR1[255:128] < binop_inR1[127:0]};
  assign main_x2_in = zll_main_dev10_in[107:8];
  Main_x2  inst (main_x2_in[99:0], main_x2_out);
  assign resize_inR2 = main_x2_out;
  assign resize_inR3 = zll_main_dev10_in[7:1];
  assign binop_inR2 = {128'(resize_inR3[6:0]), 128'h00000000000000000000000000000031};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h00000000000000000000000000000064};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[6:0];
  assign binop_inR4 = {128'(resize_inR5[6:0]), 128'h00000000000000000000000000000002};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h00000000000000000000000000000064};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[6:0];
  assign binop_inR6 = {128'(resize_inR7[6:0]), 128'h00000000000000000000000000000001};
  assign binop_inR7 = {binop_inR6[255:128] + binop_inR6[127:0], 128'h00000000000000000000000000000064};
  assign resize_inR8 = binop_inR7[255:128] % binop_inR7[127:0];
  assign resize_inR9 = resize_inR8[6:0];
  assign binop_inR8 = {128'h00000000000000000000000000000064, 128'(resize_inR9[6:0])};
  assign binop_inR9 = {binop_inR8[255:128] - binop_inR8[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR10 = {binop_inR9[255:128] - binop_inR9[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR11 = {128'(resize_inR2[99:0]), binop_inR10[255:128] * binop_inR10[127:0]};
  assign resize_inR10 = binop_inR11[255:128] >> binop_inR11[127:0];
  assign zll_main_dev9_in = {arg0, arg1, binop_in[255:128] < binop_in[127:0]};
  assign resize_inR11 = zll_main_dev9_in[107:8];
  assign resize_inR12 = zll_main_dev9_in[7:1];
  assign binop_inR12 = {128'(resize_inR12[6:0]), 128'h00000000000000000000000000000002};
  assign binop_inR13 = {binop_inR12[255:128] * binop_inR12[127:0], 128'h00000000000000000000000000000064};
  assign resize_inR13 = binop_inR13[255:128] % binop_inR13[127:0];
  assign resize_inR14 = resize_inR13[6:0];
  assign binop_inR14 = {128'(resize_inR14[6:0]), 128'h00000000000000000000000000000001};
  assign binop_inR15 = {binop_inR14[255:128] + binop_inR14[127:0], 128'h00000000000000000000000000000064};
  assign resize_inR15 = binop_inR15[255:128] % binop_inR15[127:0];
  assign resize_inR16 = resize_inR15[6:0];
  assign binop_inR16 = {128'h00000000000000000000000000000064, 128'(resize_inR16[6:0])};
  assign binop_inR17 = {binop_inR16[255:128] - binop_inR16[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR18 = {binop_inR17[255:128] - binop_inR17[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR19 = {128'(resize_inR11[99:0]), binop_inR18[255:128] * binop_inR18[127:0]};
  assign resize_inR17 = binop_inR19[255:128] >> binop_inR19[127:0];
  assign res = (zll_main_dev9_in[0] == 1'h1) ? resize_inR17[0] : resize_inR10[0];
endmodule

module Main_x2 (input logic [99:0] arg0,
  output logic [99:0] res);
  logic [199:0] binop_in;
  assign binop_in = {arg0, 100'h0000000000000000000000002};
  assign res = binop_in[199:100] * binop_in[99:0];
endmodule

module ReWire_Prelude_not (input logic [0:0] arg0,
  output logic [0:0] res);
  logic [0:0] lit_in;
  assign lit_in = arg0;
  assign res = (lit_in[0] == 1'h1) ? 1'h0 : 1'h1;
endmodule