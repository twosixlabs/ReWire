module top_level (input logic [0:0] __in0,
  output logic [0:0] __out0);
  logic [0:0] __continue;
  assign {__continue, __out0} = 1'h1;
endmodule