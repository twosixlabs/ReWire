module top_level (input logic [7:0] __in0,
  output logic [7:0] __out0);
  logic [7:0] zll_main_loop2_in;
  logic [7:0] main_myrotr_in;
  logic [15:0] zll_main_myrotr2_in;
  logic [15:0] zll_main_myrotr_in;
  logic [15:0] binop_in;
  logic [15:0] zll_main_myrotr4_in;
  logic [15:0] binop_inR1;
  logic [15:0] binop_inR2;
  logic [15:0] binop_inR3;
  logic [15:0] binop_inR4;
  logic [7:0] main_myarithrotr_in;
  logic [15:0] zll_main_myarithrotr1_in;
  logic [15:0] zll_main_myarithrotr3_in;
  logic [15:0] binop_inR5;
  logic [15:0] zll_main_myarithrotr5_in;
  logic [15:0] binop_inR6;
  logic [15:0] binop_inR7;
  logic [15:0] binop_inR8;
  logic [15:0] binop_inR9;
  logic [8:0] zll_main_loop_in;
  logic [8:0] zll_main_loop1_in;
  logic [0:0] __padding;
  assign zll_main_loop2_in = __in0;
  assign main_myrotr_in = zll_main_loop2_in[7:0];
  assign zll_main_myrotr2_in = {main_myrotr_in[7:0], 8'h3};
  assign zll_main_myrotr_in = zll_main_myrotr2_in[15:0];
  assign binop_in = {zll_main_myrotr_in[7:0], 8'h8};
  assign zll_main_myrotr4_in = {zll_main_myrotr_in[15:8], binop_in[15:8] % binop_in[7:0]};
  assign binop_inR1 = {8'h8, zll_main_myrotr4_in[7:0]};
  assign binop_inR2 = {zll_main_myrotr4_in[15:8], binop_inR1[15:8] - binop_inR1[7:0]};
  assign binop_inR3 = {zll_main_myrotr4_in[15:8], zll_main_myrotr4_in[7:0]};
  assign binop_inR4 = {binop_inR2[15:8] << binop_inR2[7:0], binop_inR3[15:8] >> binop_inR3[7:0]};
  assign main_myarithrotr_in = binop_inR4[15:8] | binop_inR4[7:0];
  assign zll_main_myarithrotr1_in = {main_myarithrotr_in[7:0], 8'h5};
  assign zll_main_myarithrotr3_in = zll_main_myarithrotr1_in[15:0];
  assign binop_inR5 = {zll_main_myarithrotr3_in[7:0], 8'h8};
  assign zll_main_myarithrotr5_in = {zll_main_myarithrotr3_in[15:8], binop_inR5[15:8] % binop_inR5[7:0]};
  assign binop_inR6 = {8'h8, zll_main_myarithrotr5_in[7:0]};
  assign binop_inR7 = {zll_main_myarithrotr5_in[15:8], binop_inR6[15:8] - binop_inR6[7:0]};
  assign binop_inR8 = {zll_main_myarithrotr5_in[15:8], zll_main_myarithrotr5_in[7:0]};
  assign binop_inR9 = {binop_inR7[15:8] << binop_inR7[7:0], binop_inR8[15:8] >>> binop_inR8[7:0]};
  assign zll_main_loop_in = {1'h0, binop_inR9[15:8] | binop_inR9[7:0]};
  assign zll_main_loop1_in = zll_main_loop_in[8:0];
  assign {__padding, __out0} = {1'h1, zll_main_loop1_in[7:0]};
endmodule