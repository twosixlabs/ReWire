module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [99:0] __in0,
  output logic [99:0] __out0);
  logic [2099:0] zll_pure_dispatch1_in;
  logic [2099:0] zll_main_dev3_in;
  logic [1099:0] main_ss$_in;
  logic [1099:0] zll_main_ss$_in;
  logic [1099:0] zll_main_ss$5_in;
  logic [999:0] id_in;
  logic [999:0] zll_main_ss$3_in;
  logic [999:0] zll_main_ss$3_out;
  logic [999:0] id_inR1;
  logic [99:0] zll_main_x2_in;
  logic [99:0] zll_main_x2_out;
  logic [999:0] id_inR2;
  logic [999:0] zll_main_ss$3_inR1;
  logic [999:0] zll_main_ss$3_outR1;
  logic [999:0] id_inR3;
  logic [99:0] zll_main_x2_inR1;
  logic [99:0] zll_main_x2_outR1;
  logic [999:0] id_inR4;
  logic [999:0] zll_main_ss$3_inR2;
  logic [999:0] zll_main_ss$3_outR2;
  logic [999:0] id_inR5;
  logic [99:0] zll_main_x2_inR2;
  logic [99:0] zll_main_x2_outR2;
  logic [999:0] id_inR6;
  logic [999:0] zll_main_ss$3_inR3;
  logic [999:0] zll_main_ss$3_outR3;
  logic [999:0] id_inR7;
  logic [99:0] zll_main_x2_inR3;
  logic [99:0] zll_main_x2_outR3;
  logic [999:0] id_inR8;
  logic [999:0] zll_main_ss$3_inR4;
  logic [999:0] zll_main_ss$3_outR4;
  logic [999:0] id_inR9;
  logic [99:0] zll_main_x2_inR4;
  logic [99:0] zll_main_x2_outR4;
  logic [999:0] id_inR10;
  logic [999:0] zll_main_ss$3_inR5;
  logic [999:0] zll_main_ss$3_outR5;
  logic [999:0] id_inR11;
  logic [99:0] zll_main_x2_inR5;
  logic [99:0] zll_main_x2_outR5;
  logic [999:0] id_inR12;
  logic [999:0] zll_main_ss$3_inR6;
  logic [999:0] zll_main_ss$3_outR6;
  logic [999:0] id_inR13;
  logic [99:0] zll_main_x2_inR6;
  logic [99:0] zll_main_x2_outR6;
  logic [999:0] id_inR14;
  logic [999:0] zll_main_ss$3_inR7;
  logic [999:0] zll_main_ss$3_outR7;
  logic [999:0] id_inR15;
  logic [99:0] zll_main_x2_inR7;
  logic [99:0] zll_main_x2_outR7;
  logic [999:0] id_inR16;
  logic [999:0] zll_main_ss$3_inR8;
  logic [999:0] zll_main_ss$3_outR8;
  logic [999:0] id_inR17;
  logic [99:0] zll_main_x2_inR8;
  logic [99:0] zll_main_x2_outR8;
  logic [999:0] id_inR18;
  logic [999:0] zll_main_ss$3_inR9;
  logic [999:0] zll_main_ss$3_outR9;
  logic [999:0] id_inR19;
  logic [99:0] zll_main_x2_inR9;
  logic [99:0] zll_main_x2_outR9;
  logic [999:0] zll_main_dev7_in;
  logic [2100:0] zll_main_dev_in;
  logic [2100:0] zll_main_dev11_in;
  logic [999:0] main_dev_in;
  logic [1999:0] zll_main_dev14_in;
  logic [1999:0] zll_main_dev10_in;
  logic [2100:0] zll_main_dev1_in;
  logic [2100:0] zll_main_dev16_in;
  logic [1999:0] zll_main_dev6_in;
  logic [999:0] zll_main_dev5_in;
  logic [999:0] id_inR20;
  logic [0:0] __continue;
  logic [999:0] __resumption_tag;
  logic [999:0] __st0;
  logic [999:0] __resumption_tag_next;
  logic [999:0] __st0_next;
  assign zll_pure_dispatch1_in = {__in0, {__resumption_tag, __st0}};
  assign zll_main_dev3_in = {zll_pure_dispatch1_in[1999:1000], zll_pure_dispatch1_in[2099:2000], zll_pure_dispatch1_in[999:0]};
  assign main_ss$_in = {zll_main_dev3_in[2099:1100], zll_main_dev3_in[1099:1000]};
  assign zll_main_ss$_in = {main_ss$_in[1099:100], main_ss$_in[99:0]};
  assign zll_main_ss$5_in = zll_main_ss$_in[1099:0];
  assign id_in = zll_main_ss$5_in[1099:100];
  assign zll_main_ss$3_in = {id_in[899:0], zll_main_ss$5_in[99:0]};
  ZLL_Main_ss$3  inst (zll_main_ss$3_in[999:100], zll_main_ss$3_in[99:0], zll_main_ss$3_out);
  assign id_inR1 = zll_main_ss$3_out;
  assign zll_main_x2_in = id_inR1[999:900];
  ZLL_Main_x2  instR1 (zll_main_x2_in[99:0], zll_main_x2_out);
  assign id_inR2 = zll_main_ss$5_in[1099:100];
  assign zll_main_ss$3_inR1 = {id_inR2[899:0], zll_main_ss$5_in[99:0]};
  ZLL_Main_ss$3  instR2 (zll_main_ss$3_inR1[999:100], zll_main_ss$3_inR1[99:0], zll_main_ss$3_outR1);
  assign id_inR3 = zll_main_ss$3_outR1;
  assign zll_main_x2_inR1 = id_inR3[899:800];
  ZLL_Main_x2  instR3 (zll_main_x2_inR1[99:0], zll_main_x2_outR1);
  assign id_inR4 = zll_main_ss$5_in[1099:100];
  assign zll_main_ss$3_inR2 = {id_inR4[899:0], zll_main_ss$5_in[99:0]};
  ZLL_Main_ss$3  instR4 (zll_main_ss$3_inR2[999:100], zll_main_ss$3_inR2[99:0], zll_main_ss$3_outR2);
  assign id_inR5 = zll_main_ss$3_outR2;
  assign zll_main_x2_inR2 = id_inR5[799:700];
  ZLL_Main_x2  instR5 (zll_main_x2_inR2[99:0], zll_main_x2_outR2);
  assign id_inR6 = zll_main_ss$5_in[1099:100];
  assign zll_main_ss$3_inR3 = {id_inR6[899:0], zll_main_ss$5_in[99:0]};
  ZLL_Main_ss$3  instR6 (zll_main_ss$3_inR3[999:100], zll_main_ss$3_inR3[99:0], zll_main_ss$3_outR3);
  assign id_inR7 = zll_main_ss$3_outR3;
  assign zll_main_x2_inR3 = id_inR7[699:600];
  ZLL_Main_x2  instR7 (zll_main_x2_inR3[99:0], zll_main_x2_outR3);
  assign id_inR8 = zll_main_ss$5_in[1099:100];
  assign zll_main_ss$3_inR4 = {id_inR8[899:0], zll_main_ss$5_in[99:0]};
  ZLL_Main_ss$3  instR8 (zll_main_ss$3_inR4[999:100], zll_main_ss$3_inR4[99:0], zll_main_ss$3_outR4);
  assign id_inR9 = zll_main_ss$3_outR4;
  assign zll_main_x2_inR4 = id_inR9[599:500];
  ZLL_Main_x2  instR9 (zll_main_x2_inR4[99:0], zll_main_x2_outR4);
  assign id_inR10 = zll_main_ss$5_in[1099:100];
  assign zll_main_ss$3_inR5 = {id_inR10[899:0], zll_main_ss$5_in[99:0]};
  ZLL_Main_ss$3  instR10 (zll_main_ss$3_inR5[999:100], zll_main_ss$3_inR5[99:0], zll_main_ss$3_outR5);
  assign id_inR11 = zll_main_ss$3_outR5;
  assign zll_main_x2_inR5 = id_inR11[499:400];
  ZLL_Main_x2  instR11 (zll_main_x2_inR5[99:0], zll_main_x2_outR5);
  assign id_inR12 = zll_main_ss$5_in[1099:100];
  assign zll_main_ss$3_inR6 = {id_inR12[899:0], zll_main_ss$5_in[99:0]};
  ZLL_Main_ss$3  instR12 (zll_main_ss$3_inR6[999:100], zll_main_ss$3_inR6[99:0], zll_main_ss$3_outR6);
  assign id_inR13 = zll_main_ss$3_outR6;
  assign zll_main_x2_inR6 = id_inR13[399:300];
  ZLL_Main_x2  instR13 (zll_main_x2_inR6[99:0], zll_main_x2_outR6);
  assign id_inR14 = zll_main_ss$5_in[1099:100];
  assign zll_main_ss$3_inR7 = {id_inR14[899:0], zll_main_ss$5_in[99:0]};
  ZLL_Main_ss$3  instR14 (zll_main_ss$3_inR7[999:100], zll_main_ss$3_inR7[99:0], zll_main_ss$3_outR7);
  assign id_inR15 = zll_main_ss$3_outR7;
  assign zll_main_x2_inR7 = id_inR15[299:200];
  ZLL_Main_x2  instR15 (zll_main_x2_inR7[99:0], zll_main_x2_outR7);
  assign id_inR16 = zll_main_ss$5_in[1099:100];
  assign zll_main_ss$3_inR8 = {id_inR16[899:0], zll_main_ss$5_in[99:0]};
  ZLL_Main_ss$3  instR16 (zll_main_ss$3_inR8[999:100], zll_main_ss$3_inR8[99:0], zll_main_ss$3_outR8);
  assign id_inR17 = zll_main_ss$3_outR8;
  assign zll_main_x2_inR8 = id_inR17[199:100];
  ZLL_Main_x2  instR17 (zll_main_x2_inR8[99:0], zll_main_x2_outR8);
  assign id_inR18 = zll_main_ss$5_in[1099:100];
  assign zll_main_ss$3_inR9 = {id_inR18[899:0], zll_main_ss$5_in[99:0]};
  ZLL_Main_ss$3  instR18 (zll_main_ss$3_inR9[999:100], zll_main_ss$3_inR9[99:0], zll_main_ss$3_outR9);
  assign id_inR19 = zll_main_ss$3_outR9;
  assign zll_main_x2_inR9 = id_inR19[99:0];
  ZLL_Main_x2  instR19 (zll_main_x2_inR9[99:0], zll_main_x2_outR9);
  assign zll_main_dev7_in = {zll_main_x2_out, zll_main_x2_outR1, zll_main_x2_outR2, zll_main_x2_outR3, zll_main_x2_outR4, zll_main_x2_outR5, zll_main_x2_outR6, zll_main_x2_outR7, zll_main_x2_outR8, zll_main_x2_outR9};
  assign zll_main_dev_in = {{101'h1, {10'h3e8{1'h0}}}, zll_main_dev7_in[999:0]};
  assign zll_main_dev11_in = zll_main_dev_in[2100:0];
  assign main_dev_in = zll_main_dev11_in[999:0];
  assign zll_main_dev14_in = {main_dev_in[999:0], main_dev_in[999:0]};
  assign zll_main_dev10_in = zll_main_dev14_in[1999:0];
  assign zll_main_dev1_in = {{7'h65{1'h0}}, zll_main_dev10_in[1999:1000], zll_main_dev10_in[999:0]};
  assign zll_main_dev16_in = zll_main_dev1_in[2100:0];
  assign zll_main_dev6_in = {zll_main_dev16_in[1999:1000], zll_main_dev16_in[999:0]};
  assign zll_main_dev5_in = zll_main_dev6_in[1999:1000];
  assign id_inR20 = zll_main_dev5_in[999:0];
  assign {__continue, __out0, __resumption_tag_next, __st0_next} = {1'h1, id_inR20[999:900], zll_main_dev6_in[1999:1000], zll_main_dev6_in[999:0]};
  initial {__resumption_tag, __st0} <= {11'h7d0{1'h0}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      {__resumption_tag, __st0} <= {11'h7d0{1'h0}};
    end else begin
      {__resumption_tag, __st0} <= {__resumption_tag_next, __st0_next};
    end
  end
endmodule

module ZLL_Main_ss$3 (input logic [899:0] arg0,
  input logic [99:0] arg1,
  output logic [999:0] res);
  logic [999:0] zll_main_ss$2_in;
  logic [999:0] id_in;
  assign zll_main_ss$2_in = {arg0, arg1};
  assign id_in = zll_main_ss$2_in[999:0];
  assign res = {id_in[999:100], id_in[99:0]};
endmodule

module ZLL_Main_x2 (input logic [99:0] arg0,
  output logic [99:0] res);
  logic [199:0] binop_in;
  assign binop_in = {arg0, 100'h2};
  assign res = binop_in[199:100] * binop_in[99:0];
endmodule