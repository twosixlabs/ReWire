module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [63:0] __in0,
  input logic [63:0] __in1,
  output logic [63:0] __out0,
  output logic [63:0] __out1);
  logic [127:0] main_loop_in;
  logic [127:0] main_compute_in;
  logic [127:0] zll_main_compute42_in;
  logic [130:0] zll_main_compute20_in;
  logic [7:0] zll_main_compute20_out;
  logic [130:0] zll_main_compute20_inR1;
  logic [7:0] zll_main_compute20_outR1;
  logic [130:0] zll_main_compute20_inR2;
  logic [7:0] zll_main_compute20_outR2;
  logic [130:0] zll_main_compute20_inR3;
  logic [7:0] zll_main_compute20_outR3;
  logic [130:0] zll_main_compute20_inR4;
  logic [7:0] zll_main_compute20_outR4;
  logic [130:0] zll_main_compute20_inR5;
  logic [7:0] zll_main_compute20_outR5;
  logic [130:0] zll_main_compute20_inR6;
  logic [7:0] zll_main_compute20_outR6;
  logic [130:0] zll_main_compute20_inR7;
  logic [7:0] zll_main_compute20_outR7;
  logic [130:0] zll_main_compute41_in;
  logic [7:0] zll_main_compute41_out;
  logic [130:0] zll_main_compute41_inR1;
  logic [7:0] zll_main_compute41_outR1;
  logic [130:0] zll_main_compute41_inR2;
  logic [7:0] zll_main_compute41_outR2;
  logic [130:0] zll_main_compute41_inR3;
  logic [7:0] zll_main_compute41_outR3;
  logic [130:0] zll_main_compute41_inR4;
  logic [7:0] zll_main_compute41_outR4;
  logic [130:0] zll_main_compute41_inR5;
  logic [7:0] zll_main_compute41_outR5;
  logic [130:0] zll_main_compute41_inR6;
  logic [7:0] zll_main_compute41_outR6;
  logic [130:0] zll_main_compute41_inR7;
  logic [7:0] zll_main_compute41_outR7;
  logic [128:0] zll_main_loop2_in;
  logic [128:0] zll_main_loop_in;
  logic [0:0] __continue;
  logic [127:0] __resumption_tag;
  logic [127:0] __resumption_tag_next;
  assign main_loop_in = __resumption_tag;
  assign main_compute_in = main_loop_in[127:0];
  assign zll_main_compute42_in = main_compute_in[127:0];
  assign zll_main_compute20_in = {zll_main_compute42_in[127:64], zll_main_compute42_in[63:0], 3'h0};
  ZLL_Main_compute20  inst (zll_main_compute20_in[130:67], zll_main_compute20_in[66:3], zll_main_compute20_in[2:0], zll_main_compute20_out);
  assign zll_main_compute20_inR1 = {zll_main_compute42_in[127:64], zll_main_compute42_in[63:0], 3'h1};
  ZLL_Main_compute20  instR1 (zll_main_compute20_inR1[130:67], zll_main_compute20_inR1[66:3], zll_main_compute20_inR1[2:0], zll_main_compute20_outR1);
  assign zll_main_compute20_inR2 = {zll_main_compute42_in[127:64], zll_main_compute42_in[63:0], 3'h2};
  ZLL_Main_compute20  instR2 (zll_main_compute20_inR2[130:67], zll_main_compute20_inR2[66:3], zll_main_compute20_inR2[2:0], zll_main_compute20_outR2);
  assign zll_main_compute20_inR3 = {zll_main_compute42_in[127:64], zll_main_compute42_in[63:0], 3'h3};
  ZLL_Main_compute20  instR3 (zll_main_compute20_inR3[130:67], zll_main_compute20_inR3[66:3], zll_main_compute20_inR3[2:0], zll_main_compute20_outR3);
  assign zll_main_compute20_inR4 = {zll_main_compute42_in[127:64], zll_main_compute42_in[63:0], 3'h4};
  ZLL_Main_compute20  instR4 (zll_main_compute20_inR4[130:67], zll_main_compute20_inR4[66:3], zll_main_compute20_inR4[2:0], zll_main_compute20_outR4);
  assign zll_main_compute20_inR5 = {zll_main_compute42_in[127:64], zll_main_compute42_in[63:0], 3'h5};
  ZLL_Main_compute20  instR5 (zll_main_compute20_inR5[130:67], zll_main_compute20_inR5[66:3], zll_main_compute20_inR5[2:0], zll_main_compute20_outR5);
  assign zll_main_compute20_inR6 = {zll_main_compute42_in[127:64], zll_main_compute42_in[63:0], 3'h6};
  ZLL_Main_compute20  instR6 (zll_main_compute20_inR6[130:67], zll_main_compute20_inR6[66:3], zll_main_compute20_inR6[2:0], zll_main_compute20_outR6);
  assign zll_main_compute20_inR7 = {zll_main_compute42_in[127:64], zll_main_compute42_in[63:0], 3'h7};
  ZLL_Main_compute20  instR7 (zll_main_compute20_inR7[130:67], zll_main_compute20_inR7[66:3], zll_main_compute20_inR7[2:0], zll_main_compute20_outR7);
  assign zll_main_compute41_in = {zll_main_compute42_in[127:64], zll_main_compute42_in[63:0], 3'h0};
  ZLL_Main_compute41  instR8 (zll_main_compute41_in[130:67], zll_main_compute41_in[66:3], zll_main_compute41_in[2:0], zll_main_compute41_out);
  assign zll_main_compute41_inR1 = {zll_main_compute42_in[127:64], zll_main_compute42_in[63:0], 3'h1};
  ZLL_Main_compute41  instR9 (zll_main_compute41_inR1[130:67], zll_main_compute41_inR1[66:3], zll_main_compute41_inR1[2:0], zll_main_compute41_outR1);
  assign zll_main_compute41_inR2 = {zll_main_compute42_in[127:64], zll_main_compute42_in[63:0], 3'h2};
  ZLL_Main_compute41  instR10 (zll_main_compute41_inR2[130:67], zll_main_compute41_inR2[66:3], zll_main_compute41_inR2[2:0], zll_main_compute41_outR2);
  assign zll_main_compute41_inR3 = {zll_main_compute42_in[127:64], zll_main_compute42_in[63:0], 3'h3};
  ZLL_Main_compute41  instR11 (zll_main_compute41_inR3[130:67], zll_main_compute41_inR3[66:3], zll_main_compute41_inR3[2:0], zll_main_compute41_outR3);
  assign zll_main_compute41_inR4 = {zll_main_compute42_in[127:64], zll_main_compute42_in[63:0], 3'h4};
  ZLL_Main_compute41  instR12 (zll_main_compute41_inR4[130:67], zll_main_compute41_inR4[66:3], zll_main_compute41_inR4[2:0], zll_main_compute41_outR4);
  assign zll_main_compute41_inR5 = {zll_main_compute42_in[127:64], zll_main_compute42_in[63:0], 3'h5};
  ZLL_Main_compute41  instR13 (zll_main_compute41_inR5[130:67], zll_main_compute41_inR5[66:3], zll_main_compute41_inR5[2:0], zll_main_compute41_outR5);
  assign zll_main_compute41_inR6 = {zll_main_compute42_in[127:64], zll_main_compute42_in[63:0], 3'h6};
  ZLL_Main_compute41  instR14 (zll_main_compute41_inR6[130:67], zll_main_compute41_inR6[66:3], zll_main_compute41_inR6[2:0], zll_main_compute41_outR6);
  assign zll_main_compute41_inR7 = {zll_main_compute42_in[127:64], zll_main_compute42_in[63:0], 3'h7};
  ZLL_Main_compute41  instR15 (zll_main_compute41_inR7[130:67], zll_main_compute41_inR7[66:3], zll_main_compute41_inR7[2:0], zll_main_compute41_outR7);
  assign zll_main_loop2_in = {1'h0, {zll_main_compute20_out, zll_main_compute20_outR1, zll_main_compute20_outR2, zll_main_compute20_outR3, zll_main_compute20_outR4, zll_main_compute20_outR5, zll_main_compute20_outR6, zll_main_compute20_outR7, zll_main_compute41_out, zll_main_compute41_outR1, zll_main_compute41_outR2, zll_main_compute41_outR3, zll_main_compute41_outR4, zll_main_compute41_outR5, zll_main_compute41_outR6, zll_main_compute41_outR7}};
  assign zll_main_loop_in = zll_main_loop2_in[128:0];
  assign {__continue, __out0, __out1, __resumption_tag_next} = {1'h1, zll_main_loop_in[127:0]};
  initial __resumption_tag <= {8'h80{1'h0}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      __resumption_tag <= {8'h80{1'h0}};
    end else begin
      __resumption_tag <= __resumption_tag_next;
    end
  end
endmodule

module ZLL_Main_compute2 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [255:0] binop_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [67:0] zll_main_compute1_in;
  logic [63:0] resize_inR2;
  logic [2:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR8;
  logic [2:0] resize_inR9;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR10;
  logic [67:0] zll_main_compute_in;
  logic [63:0] resize_inR11;
  logic [2:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [127:0] resize_inR13;
  logic [2:0] resize_inR14;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR15;
  logic [2:0] resize_inR16;
  logic [255:0] binop_inR16;
  logic [255:0] binop_inR17;
  logic [255:0] binop_inR18;
  logic [255:0] binop_inR19;
  logic [127:0] resize_inR17;
  assign resize_in = arg2;
  assign binop_in = {128'(resize_in[2:0]), 128'h00000000000000000000000000000003};
  assign resize_inR1 = arg2;
  assign binop_inR1 = {128'(resize_inR1[2:0]), 128'h00000000000000000000000000000003};
  assign zll_main_compute1_in = {arg1, arg2, binop_inR1[255:128] < binop_inR1[127:0]};
  assign resize_inR2 = zll_main_compute1_in[67:4];
  assign resize_inR3 = zll_main_compute1_in[3:1];
  assign binop_inR2 = {128'(resize_inR3[2:0]), 128'h00000000000000000000000000000003};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[2:0];
  assign binop_inR4 = {128'(resize_inR5[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR6 = {128'(resize_inR7[2:0]), 128'h00000000000000000000000000000001};
  assign binop_inR7 = {binop_inR6[255:128] + binop_inR6[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR8 = binop_inR7[255:128] % binop_inR7[127:0];
  assign resize_inR9 = resize_inR8[2:0];
  assign binop_inR8 = {128'h00000000000000000000000000000008, 128'(resize_inR9[2:0])};
  assign binop_inR9 = {binop_inR8[255:128] - binop_inR8[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR10 = {binop_inR9[255:128] - binop_inR9[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR11 = {128'(resize_inR2[63:0]), binop_inR10[255:128] * binop_inR10[127:0]};
  assign resize_inR10 = binop_inR11[255:128] >> binop_inR11[127:0];
  assign zll_main_compute_in = {arg0, arg2, binop_in[255:128] < binop_in[127:0]};
  assign resize_inR11 = zll_main_compute_in[67:4];
  assign resize_inR12 = zll_main_compute_in[3:1];
  assign binop_inR12 = {128'(resize_inR12[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR13 = {binop_inR12[255:128] * binop_inR12[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR13 = binop_inR13[255:128] % binop_inR13[127:0];
  assign resize_inR14 = resize_inR13[2:0];
  assign binop_inR14 = {128'(resize_inR14[2:0]), 128'h00000000000000000000000000000001};
  assign binop_inR15 = {binop_inR14[255:128] + binop_inR14[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR15 = binop_inR15[255:128] % binop_inR15[127:0];
  assign resize_inR16 = resize_inR15[2:0];
  assign binop_inR16 = {128'h00000000000000000000000000000008, 128'(resize_inR16[2:0])};
  assign binop_inR17 = {binop_inR16[255:128] - binop_inR16[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR18 = {binop_inR17[255:128] - binop_inR17[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR19 = {128'(resize_inR11[63:0]), binop_inR18[255:128] * binop_inR18[127:0]};
  assign resize_inR17 = binop_inR19[255:128] >> binop_inR19[127:0];
  assign res = (zll_main_compute_in[0] == 1'h1) ? resize_inR17[7:0] : resize_inR10[7:0];
endmodule

module ZLL_Main_compute6 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [255:0] binop_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [67:0] zll_main_compute5_in;
  logic [63:0] resize_inR2;
  logic [2:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR8;
  logic [67:0] zll_main_compute4_in;
  logic [63:0] resize_inR9;
  logic [2:0] resize_inR10;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR11;
  logic [2:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR13;
  assign resize_in = arg2;
  assign binop_in = {128'(resize_in[2:0]), 128'h00000000000000000000000000000003};
  assign resize_inR1 = arg2;
  assign binop_inR1 = {128'(resize_inR1[2:0]), 128'h00000000000000000000000000000003};
  assign zll_main_compute5_in = {arg2, arg1, binop_inR1[255:128] < binop_inR1[127:0]};
  assign resize_inR2 = zll_main_compute5_in[64:1];
  assign resize_inR3 = zll_main_compute5_in[67:65];
  assign binop_inR2 = {128'(resize_inR3[2:0]), 128'h00000000000000000000000000000003};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[2:0];
  assign binop_inR4 = {128'(resize_inR5[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR6 = {128'h00000000000000000000000000000008, 128'(resize_inR7[2:0])};
  assign binop_inR7 = {binop_inR6[255:128] - binop_inR6[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR8 = {binop_inR7[255:128] - binop_inR7[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR9 = {128'(resize_inR2[63:0]), binop_inR8[255:128] * binop_inR8[127:0]};
  assign resize_inR8 = binop_inR9[255:128] >> binop_inR9[127:0];
  assign zll_main_compute4_in = {arg2, arg0, binop_in[255:128] < binop_in[127:0]};
  assign resize_inR9 = zll_main_compute4_in[64:1];
  assign resize_inR10 = zll_main_compute4_in[67:65];
  assign binop_inR10 = {128'(resize_inR10[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR11 = {binop_inR10[255:128] * binop_inR10[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR11 = binop_inR11[255:128] % binop_inR11[127:0];
  assign resize_inR12 = resize_inR11[2:0];
  assign binop_inR12 = {128'h00000000000000000000000000000008, 128'(resize_inR12[2:0])};
  assign binop_inR13 = {binop_inR12[255:128] - binop_inR12[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR14 = {binop_inR13[255:128] - binop_inR13[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR15 = {128'(resize_inR9[63:0]), binop_inR14[255:128] * binop_inR14[127:0]};
  assign resize_inR13 = binop_inR15[255:128] >> binop_inR15[127:0];
  assign res = (zll_main_compute4_in[0] == 1'h1) ? resize_inR13[7:0] : resize_inR8[7:0];
endmodule

module ZLL_Main_compute8 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [255:0] binop_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [131:0] zll_main_compute7_in;
  logic [130:0] zll_main_compute6_in;
  logic [7:0] zll_main_compute6_out;
  logic [130:0] zll_main_compute6_inR1;
  logic [7:0] zll_main_compute6_outR1;
  logic [130:0] zll_main_compute6_inR2;
  logic [7:0] zll_main_compute6_outR2;
  logic [130:0] zll_main_compute6_inR3;
  logic [7:0] zll_main_compute6_outR3;
  logic [130:0] zll_main_compute6_inR4;
  logic [7:0] zll_main_compute6_outR4;
  logic [130:0] zll_main_compute6_inR5;
  logic [7:0] zll_main_compute6_outR5;
  logic [130:0] zll_main_compute6_inR6;
  logic [7:0] zll_main_compute6_outR6;
  logic [130:0] zll_main_compute6_inR7;
  logic [7:0] zll_main_compute6_outR7;
  logic [63:0] resize_inR2;
  logic [2:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR8;
  logic [131:0] zll_main_compute3_in;
  logic [130:0] zll_main_compute2_in;
  logic [7:0] zll_main_compute2_out;
  logic [130:0] zll_main_compute2_inR1;
  logic [7:0] zll_main_compute2_outR1;
  logic [130:0] zll_main_compute2_inR2;
  logic [7:0] zll_main_compute2_outR2;
  logic [130:0] zll_main_compute2_inR3;
  logic [7:0] zll_main_compute2_outR3;
  logic [130:0] zll_main_compute2_inR4;
  logic [7:0] zll_main_compute2_outR4;
  logic [130:0] zll_main_compute2_inR5;
  logic [7:0] zll_main_compute2_outR5;
  logic [130:0] zll_main_compute2_inR6;
  logic [7:0] zll_main_compute2_outR6;
  logic [130:0] zll_main_compute2_inR7;
  logic [7:0] zll_main_compute2_outR7;
  logic [63:0] resize_inR9;
  logic [2:0] resize_inR10;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR11;
  logic [2:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR13;
  assign resize_in = arg2;
  assign binop_in = {128'(resize_in[2:0]), 128'h00000000000000000000000000000003};
  assign resize_inR1 = arg2;
  assign binop_inR1 = {128'(resize_inR1[2:0]), 128'h00000000000000000000000000000003};
  assign zll_main_compute7_in = {arg0, arg1, arg2, binop_inR1[255:128] < binop_inR1[127:0]};
  assign zll_main_compute6_in = {zll_main_compute7_in[131:68], zll_main_compute7_in[67:4], 3'h0};
  ZLL_Main_compute6  inst (zll_main_compute6_in[130:67], zll_main_compute6_in[66:3], zll_main_compute6_in[2:0], zll_main_compute6_out);
  assign zll_main_compute6_inR1 = {zll_main_compute7_in[131:68], zll_main_compute7_in[67:4], 3'h1};
  ZLL_Main_compute6  instR1 (zll_main_compute6_inR1[130:67], zll_main_compute6_inR1[66:3], zll_main_compute6_inR1[2:0], zll_main_compute6_outR1);
  assign zll_main_compute6_inR2 = {zll_main_compute7_in[131:68], zll_main_compute7_in[67:4], 3'h2};
  ZLL_Main_compute6  instR2 (zll_main_compute6_inR2[130:67], zll_main_compute6_inR2[66:3], zll_main_compute6_inR2[2:0], zll_main_compute6_outR2);
  assign zll_main_compute6_inR3 = {zll_main_compute7_in[131:68], zll_main_compute7_in[67:4], 3'h3};
  ZLL_Main_compute6  instR3 (zll_main_compute6_inR3[130:67], zll_main_compute6_inR3[66:3], zll_main_compute6_inR3[2:0], zll_main_compute6_outR3);
  assign zll_main_compute6_inR4 = {zll_main_compute7_in[131:68], zll_main_compute7_in[67:4], 3'h4};
  ZLL_Main_compute6  instR4 (zll_main_compute6_inR4[130:67], zll_main_compute6_inR4[66:3], zll_main_compute6_inR4[2:0], zll_main_compute6_outR4);
  assign zll_main_compute6_inR5 = {zll_main_compute7_in[131:68], zll_main_compute7_in[67:4], 3'h5};
  ZLL_Main_compute6  instR5 (zll_main_compute6_inR5[130:67], zll_main_compute6_inR5[66:3], zll_main_compute6_inR5[2:0], zll_main_compute6_outR5);
  assign zll_main_compute6_inR6 = {zll_main_compute7_in[131:68], zll_main_compute7_in[67:4], 3'h6};
  ZLL_Main_compute6  instR6 (zll_main_compute6_inR6[130:67], zll_main_compute6_inR6[66:3], zll_main_compute6_inR6[2:0], zll_main_compute6_outR6);
  assign zll_main_compute6_inR7 = {zll_main_compute7_in[131:68], zll_main_compute7_in[67:4], 3'h7};
  ZLL_Main_compute6  instR7 (zll_main_compute6_inR7[130:67], zll_main_compute6_inR7[66:3], zll_main_compute6_inR7[2:0], zll_main_compute6_outR7);
  assign resize_inR2 = {zll_main_compute6_out, zll_main_compute6_outR1, zll_main_compute6_outR2, zll_main_compute6_outR3, zll_main_compute6_outR4, zll_main_compute6_outR5, zll_main_compute6_outR6, zll_main_compute6_outR7};
  assign resize_inR3 = zll_main_compute7_in[3:1];
  assign binop_inR2 = {128'(resize_inR3[2:0]), 128'h00000000000000000000000000000003};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[2:0];
  assign binop_inR4 = {128'(resize_inR5[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR6 = {128'h00000000000000000000000000000008, 128'(resize_inR7[2:0])};
  assign binop_inR7 = {binop_inR6[255:128] - binop_inR6[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR8 = {binop_inR7[255:128] - binop_inR7[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR9 = {128'(resize_inR2[63:0]), binop_inR8[255:128] * binop_inR8[127:0]};
  assign resize_inR8 = binop_inR9[255:128] >> binop_inR9[127:0];
  assign zll_main_compute3_in = {arg0, arg1, arg2, binop_in[255:128] < binop_in[127:0]};
  assign zll_main_compute2_in = {zll_main_compute3_in[131:68], zll_main_compute3_in[67:4], 3'h0};
  ZLL_Main_compute2  instR8 (zll_main_compute2_in[130:67], zll_main_compute2_in[66:3], zll_main_compute2_in[2:0], zll_main_compute2_out);
  assign zll_main_compute2_inR1 = {zll_main_compute3_in[131:68], zll_main_compute3_in[67:4], 3'h1};
  ZLL_Main_compute2  instR9 (zll_main_compute2_inR1[130:67], zll_main_compute2_inR1[66:3], zll_main_compute2_inR1[2:0], zll_main_compute2_outR1);
  assign zll_main_compute2_inR2 = {zll_main_compute3_in[131:68], zll_main_compute3_in[67:4], 3'h2};
  ZLL_Main_compute2  instR10 (zll_main_compute2_inR2[130:67], zll_main_compute2_inR2[66:3], zll_main_compute2_inR2[2:0], zll_main_compute2_outR2);
  assign zll_main_compute2_inR3 = {zll_main_compute3_in[131:68], zll_main_compute3_in[67:4], 3'h3};
  ZLL_Main_compute2  instR11 (zll_main_compute2_inR3[130:67], zll_main_compute2_inR3[66:3], zll_main_compute2_inR3[2:0], zll_main_compute2_outR3);
  assign zll_main_compute2_inR4 = {zll_main_compute3_in[131:68], zll_main_compute3_in[67:4], 3'h4};
  ZLL_Main_compute2  instR12 (zll_main_compute2_inR4[130:67], zll_main_compute2_inR4[66:3], zll_main_compute2_inR4[2:0], zll_main_compute2_outR4);
  assign zll_main_compute2_inR5 = {zll_main_compute3_in[131:68], zll_main_compute3_in[67:4], 3'h5};
  ZLL_Main_compute2  instR13 (zll_main_compute2_inR5[130:67], zll_main_compute2_inR5[66:3], zll_main_compute2_inR5[2:0], zll_main_compute2_outR5);
  assign zll_main_compute2_inR6 = {zll_main_compute3_in[131:68], zll_main_compute3_in[67:4], 3'h6};
  ZLL_Main_compute2  instR14 (zll_main_compute2_inR6[130:67], zll_main_compute2_inR6[66:3], zll_main_compute2_inR6[2:0], zll_main_compute2_outR6);
  assign zll_main_compute2_inR7 = {zll_main_compute3_in[131:68], zll_main_compute3_in[67:4], 3'h7};
  ZLL_Main_compute2  instR15 (zll_main_compute2_inR7[130:67], zll_main_compute2_inR7[66:3], zll_main_compute2_inR7[2:0], zll_main_compute2_outR7);
  assign resize_inR9 = {zll_main_compute2_out, zll_main_compute2_outR1, zll_main_compute2_outR2, zll_main_compute2_outR3, zll_main_compute2_outR4, zll_main_compute2_outR5, zll_main_compute2_outR6, zll_main_compute2_outR7};
  assign resize_inR10 = zll_main_compute3_in[3:1];
  assign binop_inR10 = {128'(resize_inR10[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR11 = {binop_inR10[255:128] * binop_inR10[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR11 = binop_inR11[255:128] % binop_inR11[127:0];
  assign resize_inR12 = resize_inR11[2:0];
  assign binop_inR12 = {128'h00000000000000000000000000000008, 128'(resize_inR12[2:0])};
  assign binop_inR13 = {binop_inR12[255:128] - binop_inR12[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR14 = {binop_inR13[255:128] - binop_inR13[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR15 = {128'(resize_inR9[63:0]), binop_inR14[255:128] * binop_inR14[127:0]};
  assign resize_inR13 = binop_inR15[255:128] >> binop_inR15[127:0];
  assign res = (zll_main_compute3_in[0] == 1'h1) ? resize_inR13[7:0] : resize_inR8[7:0];
endmodule

module ZLL_Main_compute16 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [255:0] binop_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [67:0] zll_main_compute15_in;
  logic [63:0] resize_inR2;
  logic [2:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR8;
  logic [67:0] zll_main_compute14_in;
  logic [63:0] resize_inR9;
  logic [2:0] resize_inR10;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR11;
  logic [2:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR13;
  assign resize_in = arg2;
  assign binop_in = {128'(resize_in[2:0]), 128'h00000000000000000000000000000003};
  assign resize_inR1 = arg2;
  assign binop_inR1 = {128'(resize_inR1[2:0]), 128'h00000000000000000000000000000003};
  assign zll_main_compute15_in = {arg1, arg2, binop_inR1[255:128] < binop_inR1[127:0]};
  assign resize_inR2 = zll_main_compute15_in[67:4];
  assign resize_inR3 = zll_main_compute15_in[3:1];
  assign binop_inR2 = {128'(resize_inR3[2:0]), 128'h00000000000000000000000000000003};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[2:0];
  assign binop_inR4 = {128'(resize_inR5[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR6 = {128'h00000000000000000000000000000008, 128'(resize_inR7[2:0])};
  assign binop_inR7 = {binop_inR6[255:128] - binop_inR6[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR8 = {binop_inR7[255:128] - binop_inR7[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR9 = {128'(resize_inR2[63:0]), binop_inR8[255:128] * binop_inR8[127:0]};
  assign resize_inR8 = binop_inR9[255:128] >> binop_inR9[127:0];
  assign zll_main_compute14_in = {arg0, arg2, binop_in[255:128] < binop_in[127:0]};
  assign resize_inR9 = zll_main_compute14_in[67:4];
  assign resize_inR10 = zll_main_compute14_in[3:1];
  assign binop_inR10 = {128'(resize_inR10[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR11 = {binop_inR10[255:128] * binop_inR10[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR11 = binop_inR11[255:128] % binop_inR11[127:0];
  assign resize_inR12 = resize_inR11[2:0];
  assign binop_inR12 = {128'h00000000000000000000000000000008, 128'(resize_inR12[2:0])};
  assign binop_inR13 = {binop_inR12[255:128] - binop_inR12[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR14 = {binop_inR13[255:128] - binop_inR13[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR15 = {128'(resize_inR9[63:0]), binop_inR14[255:128] * binop_inR14[127:0]};
  assign resize_inR13 = binop_inR15[255:128] >> binop_inR15[127:0];
  assign res = (zll_main_compute14_in[0] == 1'h1) ? resize_inR13[7:0] : resize_inR8[7:0];
endmodule

module ZLL_Main_compute18 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [255:0] binop_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [131:0] zll_main_compute17_in;
  logic [130:0] zll_main_compute16_in;
  logic [7:0] zll_main_compute16_out;
  logic [130:0] zll_main_compute16_inR1;
  logic [7:0] zll_main_compute16_outR1;
  logic [130:0] zll_main_compute16_inR2;
  logic [7:0] zll_main_compute16_outR2;
  logic [130:0] zll_main_compute16_inR3;
  logic [7:0] zll_main_compute16_outR3;
  logic [130:0] zll_main_compute16_inR4;
  logic [7:0] zll_main_compute16_outR4;
  logic [130:0] zll_main_compute16_inR5;
  logic [7:0] zll_main_compute16_outR5;
  logic [130:0] zll_main_compute16_inR6;
  logic [7:0] zll_main_compute16_outR6;
  logic [130:0] zll_main_compute16_inR7;
  logic [7:0] zll_main_compute16_outR7;
  logic [63:0] resize_inR2;
  logic [2:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR8;
  logic [2:0] resize_inR9;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR10;
  logic [131:0] zll_main_compute13_in;
  logic [130:0] zll_main_compute2_in;
  logic [7:0] zll_main_compute2_out;
  logic [130:0] zll_main_compute2_inR1;
  logic [7:0] zll_main_compute2_outR1;
  logic [130:0] zll_main_compute2_inR2;
  logic [7:0] zll_main_compute2_outR2;
  logic [130:0] zll_main_compute2_inR3;
  logic [7:0] zll_main_compute2_outR3;
  logic [130:0] zll_main_compute2_inR4;
  logic [7:0] zll_main_compute2_outR4;
  logic [130:0] zll_main_compute2_inR5;
  logic [7:0] zll_main_compute2_outR5;
  logic [130:0] zll_main_compute2_inR6;
  logic [7:0] zll_main_compute2_outR6;
  logic [130:0] zll_main_compute2_inR7;
  logic [7:0] zll_main_compute2_outR7;
  logic [63:0] resize_inR11;
  logic [2:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [127:0] resize_inR13;
  logic [2:0] resize_inR14;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR15;
  logic [2:0] resize_inR16;
  logic [255:0] binop_inR16;
  logic [255:0] binop_inR17;
  logic [255:0] binop_inR18;
  logic [255:0] binop_inR19;
  logic [127:0] resize_inR17;
  assign resize_in = arg2;
  assign binop_in = {128'(resize_in[2:0]), 128'h00000000000000000000000000000003};
  assign resize_inR1 = arg2;
  assign binop_inR1 = {128'(resize_inR1[2:0]), 128'h00000000000000000000000000000003};
  assign zll_main_compute17_in = {arg0, arg1, arg2, binop_inR1[255:128] < binop_inR1[127:0]};
  assign zll_main_compute16_in = {zll_main_compute17_in[131:68], zll_main_compute17_in[67:4], 3'h0};
  ZLL_Main_compute16  inst (zll_main_compute16_in[130:67], zll_main_compute16_in[66:3], zll_main_compute16_in[2:0], zll_main_compute16_out);
  assign zll_main_compute16_inR1 = {zll_main_compute17_in[131:68], zll_main_compute17_in[67:4], 3'h1};
  ZLL_Main_compute16  instR1 (zll_main_compute16_inR1[130:67], zll_main_compute16_inR1[66:3], zll_main_compute16_inR1[2:0], zll_main_compute16_outR1);
  assign zll_main_compute16_inR2 = {zll_main_compute17_in[131:68], zll_main_compute17_in[67:4], 3'h2};
  ZLL_Main_compute16  instR2 (zll_main_compute16_inR2[130:67], zll_main_compute16_inR2[66:3], zll_main_compute16_inR2[2:0], zll_main_compute16_outR2);
  assign zll_main_compute16_inR3 = {zll_main_compute17_in[131:68], zll_main_compute17_in[67:4], 3'h3};
  ZLL_Main_compute16  instR3 (zll_main_compute16_inR3[130:67], zll_main_compute16_inR3[66:3], zll_main_compute16_inR3[2:0], zll_main_compute16_outR3);
  assign zll_main_compute16_inR4 = {zll_main_compute17_in[131:68], zll_main_compute17_in[67:4], 3'h4};
  ZLL_Main_compute16  instR4 (zll_main_compute16_inR4[130:67], zll_main_compute16_inR4[66:3], zll_main_compute16_inR4[2:0], zll_main_compute16_outR4);
  assign zll_main_compute16_inR5 = {zll_main_compute17_in[131:68], zll_main_compute17_in[67:4], 3'h5};
  ZLL_Main_compute16  instR5 (zll_main_compute16_inR5[130:67], zll_main_compute16_inR5[66:3], zll_main_compute16_inR5[2:0], zll_main_compute16_outR5);
  assign zll_main_compute16_inR6 = {zll_main_compute17_in[131:68], zll_main_compute17_in[67:4], 3'h6};
  ZLL_Main_compute16  instR6 (zll_main_compute16_inR6[130:67], zll_main_compute16_inR6[66:3], zll_main_compute16_inR6[2:0], zll_main_compute16_outR6);
  assign zll_main_compute16_inR7 = {zll_main_compute17_in[131:68], zll_main_compute17_in[67:4], 3'h7};
  ZLL_Main_compute16  instR7 (zll_main_compute16_inR7[130:67], zll_main_compute16_inR7[66:3], zll_main_compute16_inR7[2:0], zll_main_compute16_outR7);
  assign resize_inR2 = {zll_main_compute16_out, zll_main_compute16_outR1, zll_main_compute16_outR2, zll_main_compute16_outR3, zll_main_compute16_outR4, zll_main_compute16_outR5, zll_main_compute16_outR6, zll_main_compute16_outR7};
  assign resize_inR3 = zll_main_compute17_in[3:1];
  assign binop_inR2 = {128'(resize_inR3[2:0]), 128'h00000000000000000000000000000003};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[2:0];
  assign binop_inR4 = {128'(resize_inR5[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR6 = {128'(resize_inR7[2:0]), 128'h00000000000000000000000000000001};
  assign binop_inR7 = {binop_inR6[255:128] + binop_inR6[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR8 = binop_inR7[255:128] % binop_inR7[127:0];
  assign resize_inR9 = resize_inR8[2:0];
  assign binop_inR8 = {128'h00000000000000000000000000000008, 128'(resize_inR9[2:0])};
  assign binop_inR9 = {binop_inR8[255:128] - binop_inR8[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR10 = {binop_inR9[255:128] - binop_inR9[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR11 = {128'(resize_inR2[63:0]), binop_inR10[255:128] * binop_inR10[127:0]};
  assign resize_inR10 = binop_inR11[255:128] >> binop_inR11[127:0];
  assign zll_main_compute13_in = {arg0, arg1, arg2, binop_in[255:128] < binop_in[127:0]};
  assign zll_main_compute2_in = {zll_main_compute13_in[131:68], zll_main_compute13_in[67:4], 3'h0};
  ZLL_Main_compute2  instR8 (zll_main_compute2_in[130:67], zll_main_compute2_in[66:3], zll_main_compute2_in[2:0], zll_main_compute2_out);
  assign zll_main_compute2_inR1 = {zll_main_compute13_in[131:68], zll_main_compute13_in[67:4], 3'h1};
  ZLL_Main_compute2  instR9 (zll_main_compute2_inR1[130:67], zll_main_compute2_inR1[66:3], zll_main_compute2_inR1[2:0], zll_main_compute2_outR1);
  assign zll_main_compute2_inR2 = {zll_main_compute13_in[131:68], zll_main_compute13_in[67:4], 3'h2};
  ZLL_Main_compute2  instR10 (zll_main_compute2_inR2[130:67], zll_main_compute2_inR2[66:3], zll_main_compute2_inR2[2:0], zll_main_compute2_outR2);
  assign zll_main_compute2_inR3 = {zll_main_compute13_in[131:68], zll_main_compute13_in[67:4], 3'h3};
  ZLL_Main_compute2  instR11 (zll_main_compute2_inR3[130:67], zll_main_compute2_inR3[66:3], zll_main_compute2_inR3[2:0], zll_main_compute2_outR3);
  assign zll_main_compute2_inR4 = {zll_main_compute13_in[131:68], zll_main_compute13_in[67:4], 3'h4};
  ZLL_Main_compute2  instR12 (zll_main_compute2_inR4[130:67], zll_main_compute2_inR4[66:3], zll_main_compute2_inR4[2:0], zll_main_compute2_outR4);
  assign zll_main_compute2_inR5 = {zll_main_compute13_in[131:68], zll_main_compute13_in[67:4], 3'h5};
  ZLL_Main_compute2  instR13 (zll_main_compute2_inR5[130:67], zll_main_compute2_inR5[66:3], zll_main_compute2_inR5[2:0], zll_main_compute2_outR5);
  assign zll_main_compute2_inR6 = {zll_main_compute13_in[131:68], zll_main_compute13_in[67:4], 3'h6};
  ZLL_Main_compute2  instR14 (zll_main_compute2_inR6[130:67], zll_main_compute2_inR6[66:3], zll_main_compute2_inR6[2:0], zll_main_compute2_outR6);
  assign zll_main_compute2_inR7 = {zll_main_compute13_in[131:68], zll_main_compute13_in[67:4], 3'h7};
  ZLL_Main_compute2  instR15 (zll_main_compute2_inR7[130:67], zll_main_compute2_inR7[66:3], zll_main_compute2_inR7[2:0], zll_main_compute2_outR7);
  assign resize_inR11 = {zll_main_compute2_out, zll_main_compute2_outR1, zll_main_compute2_outR2, zll_main_compute2_outR3, zll_main_compute2_outR4, zll_main_compute2_outR5, zll_main_compute2_outR6, zll_main_compute2_outR7};
  assign resize_inR12 = zll_main_compute13_in[3:1];
  assign binop_inR12 = {128'(resize_inR12[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR13 = {binop_inR12[255:128] * binop_inR12[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR13 = binop_inR13[255:128] % binop_inR13[127:0];
  assign resize_inR14 = resize_inR13[2:0];
  assign binop_inR14 = {128'(resize_inR14[2:0]), 128'h00000000000000000000000000000001};
  assign binop_inR15 = {binop_inR14[255:128] + binop_inR14[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR15 = binop_inR15[255:128] % binop_inR15[127:0];
  assign resize_inR16 = resize_inR15[2:0];
  assign binop_inR16 = {128'h00000000000000000000000000000008, 128'(resize_inR16[2:0])};
  assign binop_inR17 = {binop_inR16[255:128] - binop_inR16[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR18 = {binop_inR17[255:128] - binop_inR17[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR19 = {128'(resize_inR11[63:0]), binop_inR18[255:128] * binop_inR18[127:0]};
  assign resize_inR17 = binop_inR19[255:128] >> binop_inR19[127:0];
  assign res = (zll_main_compute13_in[0] == 1'h1) ? resize_inR17[7:0] : resize_inR10[7:0];
endmodule

module ZLL_Main_compute20 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [127:0] resize_inR1;
  logic [0:0] msbit_in;
  logic [0:0] rewire_prelude_not_in;
  logic [0:0] rewire_prelude_not_out;
  logic [2:0] resize_inR2;
  logic [127:0] resize_inR3;
  logic [0:0] msbit_inR1;
  logic [0:0] rewire_prelude_not_inR1;
  logic [0:0] rewire_prelude_not_outR1;
  logic [131:0] zll_main_compute19_in;
  logic [130:0] zll_main_compute18_in;
  logic [7:0] zll_main_compute18_out;
  logic [130:0] zll_main_compute18_inR1;
  logic [7:0] zll_main_compute18_outR1;
  logic [130:0] zll_main_compute18_inR2;
  logic [7:0] zll_main_compute18_outR2;
  logic [130:0] zll_main_compute18_inR3;
  logic [7:0] zll_main_compute18_outR3;
  logic [130:0] zll_main_compute18_inR4;
  logic [7:0] zll_main_compute18_outR4;
  logic [130:0] zll_main_compute18_inR5;
  logic [7:0] zll_main_compute18_outR5;
  logic [130:0] zll_main_compute18_inR6;
  logic [7:0] zll_main_compute18_outR6;
  logic [130:0] zll_main_compute18_inR7;
  logic [7:0] zll_main_compute18_outR7;
  logic [63:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR8;
  logic [2:0] resize_inR9;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR10;
  logic [131:0] zll_main_compute9_in;
  logic [130:0] zll_main_compute8_in;
  logic [7:0] zll_main_compute8_out;
  logic [130:0] zll_main_compute8_inR1;
  logic [7:0] zll_main_compute8_outR1;
  logic [130:0] zll_main_compute8_inR2;
  logic [7:0] zll_main_compute8_outR2;
  logic [130:0] zll_main_compute8_inR3;
  logic [7:0] zll_main_compute8_outR3;
  logic [130:0] zll_main_compute8_inR4;
  logic [7:0] zll_main_compute8_outR4;
  logic [130:0] zll_main_compute8_inR5;
  logic [7:0] zll_main_compute8_outR5;
  logic [130:0] zll_main_compute8_inR6;
  logic [7:0] zll_main_compute8_outR6;
  logic [130:0] zll_main_compute8_inR7;
  logic [7:0] zll_main_compute8_outR7;
  logic [63:0] resize_inR11;
  logic [2:0] resize_inR12;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR13;
  logic [2:0] resize_inR14;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [127:0] resize_inR15;
  assign resize_in = arg2;
  assign resize_inR1 = 128'(resize_in[2:0]);
  assign msbit_in = resize_inR1[0];
  assign rewire_prelude_not_in = msbit_in[0];
  ReWire_Prelude_not  inst (rewire_prelude_not_in[0], rewire_prelude_not_out);
  assign resize_inR2 = arg2;
  assign resize_inR3 = 128'(resize_inR2[2:0]);
  assign msbit_inR1 = resize_inR3[0];
  assign rewire_prelude_not_inR1 = msbit_inR1[0];
  ReWire_Prelude_not  instR1 (rewire_prelude_not_inR1[0], rewire_prelude_not_outR1);
  assign zll_main_compute19_in = {arg0, arg1, arg2, rewire_prelude_not_outR1};
  assign zll_main_compute18_in = {zll_main_compute19_in[131:68], zll_main_compute19_in[67:4], 3'h0};
  ZLL_Main_compute18  instR2 (zll_main_compute18_in[130:67], zll_main_compute18_in[66:3], zll_main_compute18_in[2:0], zll_main_compute18_out);
  assign zll_main_compute18_inR1 = {zll_main_compute19_in[131:68], zll_main_compute19_in[67:4], 3'h1};
  ZLL_Main_compute18  instR3 (zll_main_compute18_inR1[130:67], zll_main_compute18_inR1[66:3], zll_main_compute18_inR1[2:0], zll_main_compute18_outR1);
  assign zll_main_compute18_inR2 = {zll_main_compute19_in[131:68], zll_main_compute19_in[67:4], 3'h2};
  ZLL_Main_compute18  instR4 (zll_main_compute18_inR2[130:67], zll_main_compute18_inR2[66:3], zll_main_compute18_inR2[2:0], zll_main_compute18_outR2);
  assign zll_main_compute18_inR3 = {zll_main_compute19_in[131:68], zll_main_compute19_in[67:4], 3'h3};
  ZLL_Main_compute18  instR5 (zll_main_compute18_inR3[130:67], zll_main_compute18_inR3[66:3], zll_main_compute18_inR3[2:0], zll_main_compute18_outR3);
  assign zll_main_compute18_inR4 = {zll_main_compute19_in[131:68], zll_main_compute19_in[67:4], 3'h4};
  ZLL_Main_compute18  instR6 (zll_main_compute18_inR4[130:67], zll_main_compute18_inR4[66:3], zll_main_compute18_inR4[2:0], zll_main_compute18_outR4);
  assign zll_main_compute18_inR5 = {zll_main_compute19_in[131:68], zll_main_compute19_in[67:4], 3'h5};
  ZLL_Main_compute18  instR7 (zll_main_compute18_inR5[130:67], zll_main_compute18_inR5[66:3], zll_main_compute18_inR5[2:0], zll_main_compute18_outR5);
  assign zll_main_compute18_inR6 = {zll_main_compute19_in[131:68], zll_main_compute19_in[67:4], 3'h6};
  ZLL_Main_compute18  instR8 (zll_main_compute18_inR6[130:67], zll_main_compute18_inR6[66:3], zll_main_compute18_inR6[2:0], zll_main_compute18_outR6);
  assign zll_main_compute18_inR7 = {zll_main_compute19_in[131:68], zll_main_compute19_in[67:4], 3'h7};
  ZLL_Main_compute18  instR9 (zll_main_compute18_inR7[130:67], zll_main_compute18_inR7[66:3], zll_main_compute18_inR7[2:0], zll_main_compute18_outR7);
  assign resize_inR4 = {zll_main_compute18_out, zll_main_compute18_outR1, zll_main_compute18_outR2, zll_main_compute18_outR3, zll_main_compute18_outR4, zll_main_compute18_outR5, zll_main_compute18_outR6, zll_main_compute18_outR7};
  assign resize_inR5 = zll_main_compute19_in[3:1];
  assign binop_in = {128'(resize_inR5[2:0]), 128'h00000000000000000000000000000001};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR6 = binop_inR1[255:128] % binop_inR1[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR2 = {128'(resize_inR7[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR3 = {binop_inR2[255:128] / binop_inR2[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR8 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR9 = resize_inR8[2:0];
  assign binop_inR4 = {128'h00000000000000000000000000000008, 128'(resize_inR9[2:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR7 = {128'(resize_inR4[63:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR10 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign zll_main_compute9_in = {arg0, arg1, arg2, rewire_prelude_not_out};
  assign zll_main_compute8_in = {zll_main_compute9_in[131:68], zll_main_compute9_in[67:4], 3'h0};
  ZLL_Main_compute8  instR10 (zll_main_compute8_in[130:67], zll_main_compute8_in[66:3], zll_main_compute8_in[2:0], zll_main_compute8_out);
  assign zll_main_compute8_inR1 = {zll_main_compute9_in[131:68], zll_main_compute9_in[67:4], 3'h1};
  ZLL_Main_compute8  instR11 (zll_main_compute8_inR1[130:67], zll_main_compute8_inR1[66:3], zll_main_compute8_inR1[2:0], zll_main_compute8_outR1);
  assign zll_main_compute8_inR2 = {zll_main_compute9_in[131:68], zll_main_compute9_in[67:4], 3'h2};
  ZLL_Main_compute8  instR12 (zll_main_compute8_inR2[130:67], zll_main_compute8_inR2[66:3], zll_main_compute8_inR2[2:0], zll_main_compute8_outR2);
  assign zll_main_compute8_inR3 = {zll_main_compute9_in[131:68], zll_main_compute9_in[67:4], 3'h3};
  ZLL_Main_compute8  instR13 (zll_main_compute8_inR3[130:67], zll_main_compute8_inR3[66:3], zll_main_compute8_inR3[2:0], zll_main_compute8_outR3);
  assign zll_main_compute8_inR4 = {zll_main_compute9_in[131:68], zll_main_compute9_in[67:4], 3'h4};
  ZLL_Main_compute8  instR14 (zll_main_compute8_inR4[130:67], zll_main_compute8_inR4[66:3], zll_main_compute8_inR4[2:0], zll_main_compute8_outR4);
  assign zll_main_compute8_inR5 = {zll_main_compute9_in[131:68], zll_main_compute9_in[67:4], 3'h5};
  ZLL_Main_compute8  instR15 (zll_main_compute8_inR5[130:67], zll_main_compute8_inR5[66:3], zll_main_compute8_inR5[2:0], zll_main_compute8_outR5);
  assign zll_main_compute8_inR6 = {zll_main_compute9_in[131:68], zll_main_compute9_in[67:4], 3'h6};
  ZLL_Main_compute8  instR16 (zll_main_compute8_inR6[130:67], zll_main_compute8_inR6[66:3], zll_main_compute8_inR6[2:0], zll_main_compute8_outR6);
  assign zll_main_compute8_inR7 = {zll_main_compute9_in[131:68], zll_main_compute9_in[67:4], 3'h7};
  ZLL_Main_compute8  instR17 (zll_main_compute8_inR7[130:67], zll_main_compute8_inR7[66:3], zll_main_compute8_inR7[2:0], zll_main_compute8_outR7);
  assign resize_inR11 = {zll_main_compute8_out, zll_main_compute8_outR1, zll_main_compute8_outR2, zll_main_compute8_outR3, zll_main_compute8_outR4, zll_main_compute8_outR5, zll_main_compute8_outR6, zll_main_compute8_outR7};
  assign resize_inR12 = zll_main_compute9_in[3:1];
  assign binop_inR8 = {128'(resize_inR12[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR9 = {binop_inR8[255:128] / binop_inR8[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR13 = binop_inR9[255:128] % binop_inR9[127:0];
  assign resize_inR14 = resize_inR13[2:0];
  assign binop_inR10 = {128'h00000000000000000000000000000008, 128'(resize_inR14[2:0])};
  assign binop_inR11 = {binop_inR10[255:128] - binop_inR10[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR12 = {binop_inR11[255:128] - binop_inR11[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR13 = {128'(resize_inR11[63:0]), binop_inR12[255:128] * binop_inR12[127:0]};
  assign resize_inR15 = binop_inR13[255:128] >> binop_inR13[127:0];
  assign res = (zll_main_compute9_in[0] == 1'h1) ? resize_inR15[7:0] : resize_inR10[7:0];
endmodule

module ZLL_Main_compute29 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [255:0] binop_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [131:0] zll_main_compute28_in;
  logic [130:0] zll_main_compute16_in;
  logic [7:0] zll_main_compute16_out;
  logic [130:0] zll_main_compute16_inR1;
  logic [7:0] zll_main_compute16_outR1;
  logic [130:0] zll_main_compute16_inR2;
  logic [7:0] zll_main_compute16_outR2;
  logic [130:0] zll_main_compute16_inR3;
  logic [7:0] zll_main_compute16_outR3;
  logic [130:0] zll_main_compute16_inR4;
  logic [7:0] zll_main_compute16_outR4;
  logic [130:0] zll_main_compute16_inR5;
  logic [7:0] zll_main_compute16_outR5;
  logic [130:0] zll_main_compute16_inR6;
  logic [7:0] zll_main_compute16_outR6;
  logic [130:0] zll_main_compute16_inR7;
  logic [7:0] zll_main_compute16_outR7;
  logic [63:0] resize_inR2;
  logic [2:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR8;
  logic [131:0] zll_main_compute24_in;
  logic [130:0] zll_main_compute2_in;
  logic [7:0] zll_main_compute2_out;
  logic [130:0] zll_main_compute2_inR1;
  logic [7:0] zll_main_compute2_outR1;
  logic [130:0] zll_main_compute2_inR2;
  logic [7:0] zll_main_compute2_outR2;
  logic [130:0] zll_main_compute2_inR3;
  logic [7:0] zll_main_compute2_outR3;
  logic [130:0] zll_main_compute2_inR4;
  logic [7:0] zll_main_compute2_outR4;
  logic [130:0] zll_main_compute2_inR5;
  logic [7:0] zll_main_compute2_outR5;
  logic [130:0] zll_main_compute2_inR6;
  logic [7:0] zll_main_compute2_outR6;
  logic [130:0] zll_main_compute2_inR7;
  logic [7:0] zll_main_compute2_outR7;
  logic [63:0] resize_inR9;
  logic [2:0] resize_inR10;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR11;
  logic [2:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR13;
  assign resize_in = arg2;
  assign binop_in = {128'(resize_in[2:0]), 128'h00000000000000000000000000000003};
  assign resize_inR1 = arg2;
  assign binop_inR1 = {128'(resize_inR1[2:0]), 128'h00000000000000000000000000000003};
  assign zll_main_compute28_in = {arg2, arg0, arg1, binop_inR1[255:128] < binop_inR1[127:0]};
  assign zll_main_compute16_in = {zll_main_compute28_in[128:65], zll_main_compute28_in[64:1], 3'h0};
  ZLL_Main_compute16  inst (zll_main_compute16_in[130:67], zll_main_compute16_in[66:3], zll_main_compute16_in[2:0], zll_main_compute16_out);
  assign zll_main_compute16_inR1 = {zll_main_compute28_in[128:65], zll_main_compute28_in[64:1], 3'h1};
  ZLL_Main_compute16  instR1 (zll_main_compute16_inR1[130:67], zll_main_compute16_inR1[66:3], zll_main_compute16_inR1[2:0], zll_main_compute16_outR1);
  assign zll_main_compute16_inR2 = {zll_main_compute28_in[128:65], zll_main_compute28_in[64:1], 3'h2};
  ZLL_Main_compute16  instR2 (zll_main_compute16_inR2[130:67], zll_main_compute16_inR2[66:3], zll_main_compute16_inR2[2:0], zll_main_compute16_outR2);
  assign zll_main_compute16_inR3 = {zll_main_compute28_in[128:65], zll_main_compute28_in[64:1], 3'h3};
  ZLL_Main_compute16  instR3 (zll_main_compute16_inR3[130:67], zll_main_compute16_inR3[66:3], zll_main_compute16_inR3[2:0], zll_main_compute16_outR3);
  assign zll_main_compute16_inR4 = {zll_main_compute28_in[128:65], zll_main_compute28_in[64:1], 3'h4};
  ZLL_Main_compute16  instR4 (zll_main_compute16_inR4[130:67], zll_main_compute16_inR4[66:3], zll_main_compute16_inR4[2:0], zll_main_compute16_outR4);
  assign zll_main_compute16_inR5 = {zll_main_compute28_in[128:65], zll_main_compute28_in[64:1], 3'h5};
  ZLL_Main_compute16  instR5 (zll_main_compute16_inR5[130:67], zll_main_compute16_inR5[66:3], zll_main_compute16_inR5[2:0], zll_main_compute16_outR5);
  assign zll_main_compute16_inR6 = {zll_main_compute28_in[128:65], zll_main_compute28_in[64:1], 3'h6};
  ZLL_Main_compute16  instR6 (zll_main_compute16_inR6[130:67], zll_main_compute16_inR6[66:3], zll_main_compute16_inR6[2:0], zll_main_compute16_outR6);
  assign zll_main_compute16_inR7 = {zll_main_compute28_in[128:65], zll_main_compute28_in[64:1], 3'h7};
  ZLL_Main_compute16  instR7 (zll_main_compute16_inR7[130:67], zll_main_compute16_inR7[66:3], zll_main_compute16_inR7[2:0], zll_main_compute16_outR7);
  assign resize_inR2 = {zll_main_compute16_out, zll_main_compute16_outR1, zll_main_compute16_outR2, zll_main_compute16_outR3, zll_main_compute16_outR4, zll_main_compute16_outR5, zll_main_compute16_outR6, zll_main_compute16_outR7};
  assign resize_inR3 = zll_main_compute28_in[131:129];
  assign binop_inR2 = {128'(resize_inR3[2:0]), 128'h00000000000000000000000000000003};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[2:0];
  assign binop_inR4 = {128'(resize_inR5[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR6 = {128'h00000000000000000000000000000008, 128'(resize_inR7[2:0])};
  assign binop_inR7 = {binop_inR6[255:128] - binop_inR6[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR8 = {binop_inR7[255:128] - binop_inR7[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR9 = {128'(resize_inR2[63:0]), binop_inR8[255:128] * binop_inR8[127:0]};
  assign resize_inR8 = binop_inR9[255:128] >> binop_inR9[127:0];
  assign zll_main_compute24_in = {arg2, arg0, arg1, binop_in[255:128] < binop_in[127:0]};
  assign zll_main_compute2_in = {zll_main_compute24_in[128:65], zll_main_compute24_in[64:1], 3'h0};
  ZLL_Main_compute2  instR8 (zll_main_compute2_in[130:67], zll_main_compute2_in[66:3], zll_main_compute2_in[2:0], zll_main_compute2_out);
  assign zll_main_compute2_inR1 = {zll_main_compute24_in[128:65], zll_main_compute24_in[64:1], 3'h1};
  ZLL_Main_compute2  instR9 (zll_main_compute2_inR1[130:67], zll_main_compute2_inR1[66:3], zll_main_compute2_inR1[2:0], zll_main_compute2_outR1);
  assign zll_main_compute2_inR2 = {zll_main_compute24_in[128:65], zll_main_compute24_in[64:1], 3'h2};
  ZLL_Main_compute2  instR10 (zll_main_compute2_inR2[130:67], zll_main_compute2_inR2[66:3], zll_main_compute2_inR2[2:0], zll_main_compute2_outR2);
  assign zll_main_compute2_inR3 = {zll_main_compute24_in[128:65], zll_main_compute24_in[64:1], 3'h3};
  ZLL_Main_compute2  instR11 (zll_main_compute2_inR3[130:67], zll_main_compute2_inR3[66:3], zll_main_compute2_inR3[2:0], zll_main_compute2_outR3);
  assign zll_main_compute2_inR4 = {zll_main_compute24_in[128:65], zll_main_compute24_in[64:1], 3'h4};
  ZLL_Main_compute2  instR12 (zll_main_compute2_inR4[130:67], zll_main_compute2_inR4[66:3], zll_main_compute2_inR4[2:0], zll_main_compute2_outR4);
  assign zll_main_compute2_inR5 = {zll_main_compute24_in[128:65], zll_main_compute24_in[64:1], 3'h5};
  ZLL_Main_compute2  instR13 (zll_main_compute2_inR5[130:67], zll_main_compute2_inR5[66:3], zll_main_compute2_inR5[2:0], zll_main_compute2_outR5);
  assign zll_main_compute2_inR6 = {zll_main_compute24_in[128:65], zll_main_compute24_in[64:1], 3'h6};
  ZLL_Main_compute2  instR14 (zll_main_compute2_inR6[130:67], zll_main_compute2_inR6[66:3], zll_main_compute2_inR6[2:0], zll_main_compute2_outR6);
  assign zll_main_compute2_inR7 = {zll_main_compute24_in[128:65], zll_main_compute24_in[64:1], 3'h7};
  ZLL_Main_compute2  instR15 (zll_main_compute2_inR7[130:67], zll_main_compute2_inR7[66:3], zll_main_compute2_inR7[2:0], zll_main_compute2_outR7);
  assign resize_inR9 = {zll_main_compute2_out, zll_main_compute2_outR1, zll_main_compute2_outR2, zll_main_compute2_outR3, zll_main_compute2_outR4, zll_main_compute2_outR5, zll_main_compute2_outR6, zll_main_compute2_outR7};
  assign resize_inR10 = zll_main_compute24_in[131:129];
  assign binop_inR10 = {128'(resize_inR10[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR11 = {binop_inR10[255:128] * binop_inR10[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR11 = binop_inR11[255:128] % binop_inR11[127:0];
  assign resize_inR12 = resize_inR11[2:0];
  assign binop_inR12 = {128'h00000000000000000000000000000008, 128'(resize_inR12[2:0])};
  assign binop_inR13 = {binop_inR12[255:128] - binop_inR12[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR14 = {binop_inR13[255:128] - binop_inR13[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR15 = {128'(resize_inR9[63:0]), binop_inR14[255:128] * binop_inR14[127:0]};
  assign resize_inR13 = binop_inR15[255:128] >> binop_inR15[127:0];
  assign res = (zll_main_compute24_in[0] == 1'h1) ? resize_inR13[7:0] : resize_inR8[7:0];
endmodule

module ZLL_Main_compute39 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [255:0] binop_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [131:0] zll_main_compute38_in;
  logic [130:0] zll_main_compute16_in;
  logic [7:0] zll_main_compute16_out;
  logic [130:0] zll_main_compute16_inR1;
  logic [7:0] zll_main_compute16_outR1;
  logic [130:0] zll_main_compute16_inR2;
  logic [7:0] zll_main_compute16_outR2;
  logic [130:0] zll_main_compute16_inR3;
  logic [7:0] zll_main_compute16_outR3;
  logic [130:0] zll_main_compute16_inR4;
  logic [7:0] zll_main_compute16_outR4;
  logic [130:0] zll_main_compute16_inR5;
  logic [7:0] zll_main_compute16_outR5;
  logic [130:0] zll_main_compute16_inR6;
  logic [7:0] zll_main_compute16_outR6;
  logic [130:0] zll_main_compute16_inR7;
  logic [7:0] zll_main_compute16_outR7;
  logic [63:0] resize_inR2;
  logic [2:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR8;
  logic [2:0] resize_inR9;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR10;
  logic [131:0] zll_main_compute34_in;
  logic [130:0] zll_main_compute2_in;
  logic [7:0] zll_main_compute2_out;
  logic [130:0] zll_main_compute2_inR1;
  logic [7:0] zll_main_compute2_outR1;
  logic [130:0] zll_main_compute2_inR2;
  logic [7:0] zll_main_compute2_outR2;
  logic [130:0] zll_main_compute2_inR3;
  logic [7:0] zll_main_compute2_outR3;
  logic [130:0] zll_main_compute2_inR4;
  logic [7:0] zll_main_compute2_outR4;
  logic [130:0] zll_main_compute2_inR5;
  logic [7:0] zll_main_compute2_outR5;
  logic [130:0] zll_main_compute2_inR6;
  logic [7:0] zll_main_compute2_outR6;
  logic [130:0] zll_main_compute2_inR7;
  logic [7:0] zll_main_compute2_outR7;
  logic [63:0] resize_inR11;
  logic [2:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [127:0] resize_inR13;
  logic [2:0] resize_inR14;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR15;
  logic [2:0] resize_inR16;
  logic [255:0] binop_inR16;
  logic [255:0] binop_inR17;
  logic [255:0] binop_inR18;
  logic [255:0] binop_inR19;
  logic [127:0] resize_inR17;
  assign resize_in = arg2;
  assign binop_in = {128'(resize_in[2:0]), 128'h00000000000000000000000000000003};
  assign resize_inR1 = arg2;
  assign binop_inR1 = {128'(resize_inR1[2:0]), 128'h00000000000000000000000000000003};
  assign zll_main_compute38_in = {arg2, arg0, arg1, binop_inR1[255:128] < binop_inR1[127:0]};
  assign zll_main_compute16_in = {zll_main_compute38_in[128:65], zll_main_compute38_in[64:1], 3'h0};
  ZLL_Main_compute16  inst (zll_main_compute16_in[130:67], zll_main_compute16_in[66:3], zll_main_compute16_in[2:0], zll_main_compute16_out);
  assign zll_main_compute16_inR1 = {zll_main_compute38_in[128:65], zll_main_compute38_in[64:1], 3'h1};
  ZLL_Main_compute16  instR1 (zll_main_compute16_inR1[130:67], zll_main_compute16_inR1[66:3], zll_main_compute16_inR1[2:0], zll_main_compute16_outR1);
  assign zll_main_compute16_inR2 = {zll_main_compute38_in[128:65], zll_main_compute38_in[64:1], 3'h2};
  ZLL_Main_compute16  instR2 (zll_main_compute16_inR2[130:67], zll_main_compute16_inR2[66:3], zll_main_compute16_inR2[2:0], zll_main_compute16_outR2);
  assign zll_main_compute16_inR3 = {zll_main_compute38_in[128:65], zll_main_compute38_in[64:1], 3'h3};
  ZLL_Main_compute16  instR3 (zll_main_compute16_inR3[130:67], zll_main_compute16_inR3[66:3], zll_main_compute16_inR3[2:0], zll_main_compute16_outR3);
  assign zll_main_compute16_inR4 = {zll_main_compute38_in[128:65], zll_main_compute38_in[64:1], 3'h4};
  ZLL_Main_compute16  instR4 (zll_main_compute16_inR4[130:67], zll_main_compute16_inR4[66:3], zll_main_compute16_inR4[2:0], zll_main_compute16_outR4);
  assign zll_main_compute16_inR5 = {zll_main_compute38_in[128:65], zll_main_compute38_in[64:1], 3'h5};
  ZLL_Main_compute16  instR5 (zll_main_compute16_inR5[130:67], zll_main_compute16_inR5[66:3], zll_main_compute16_inR5[2:0], zll_main_compute16_outR5);
  assign zll_main_compute16_inR6 = {zll_main_compute38_in[128:65], zll_main_compute38_in[64:1], 3'h6};
  ZLL_Main_compute16  instR6 (zll_main_compute16_inR6[130:67], zll_main_compute16_inR6[66:3], zll_main_compute16_inR6[2:0], zll_main_compute16_outR6);
  assign zll_main_compute16_inR7 = {zll_main_compute38_in[128:65], zll_main_compute38_in[64:1], 3'h7};
  ZLL_Main_compute16  instR7 (zll_main_compute16_inR7[130:67], zll_main_compute16_inR7[66:3], zll_main_compute16_inR7[2:0], zll_main_compute16_outR7);
  assign resize_inR2 = {zll_main_compute16_out, zll_main_compute16_outR1, zll_main_compute16_outR2, zll_main_compute16_outR3, zll_main_compute16_outR4, zll_main_compute16_outR5, zll_main_compute16_outR6, zll_main_compute16_outR7};
  assign resize_inR3 = zll_main_compute38_in[131:129];
  assign binop_inR2 = {128'(resize_inR3[2:0]), 128'h00000000000000000000000000000003};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[2:0];
  assign binop_inR4 = {128'(resize_inR5[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR6 = {128'(resize_inR7[2:0]), 128'h00000000000000000000000000000001};
  assign binop_inR7 = {binop_inR6[255:128] + binop_inR6[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR8 = binop_inR7[255:128] % binop_inR7[127:0];
  assign resize_inR9 = resize_inR8[2:0];
  assign binop_inR8 = {128'h00000000000000000000000000000008, 128'(resize_inR9[2:0])};
  assign binop_inR9 = {binop_inR8[255:128] - binop_inR8[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR10 = {binop_inR9[255:128] - binop_inR9[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR11 = {128'(resize_inR2[63:0]), binop_inR10[255:128] * binop_inR10[127:0]};
  assign resize_inR10 = binop_inR11[255:128] >> binop_inR11[127:0];
  assign zll_main_compute34_in = {arg2, arg0, arg1, binop_in[255:128] < binop_in[127:0]};
  assign zll_main_compute2_in = {zll_main_compute34_in[128:65], zll_main_compute34_in[64:1], 3'h0};
  ZLL_Main_compute2  instR8 (zll_main_compute2_in[130:67], zll_main_compute2_in[66:3], zll_main_compute2_in[2:0], zll_main_compute2_out);
  assign zll_main_compute2_inR1 = {zll_main_compute34_in[128:65], zll_main_compute34_in[64:1], 3'h1};
  ZLL_Main_compute2  instR9 (zll_main_compute2_inR1[130:67], zll_main_compute2_inR1[66:3], zll_main_compute2_inR1[2:0], zll_main_compute2_outR1);
  assign zll_main_compute2_inR2 = {zll_main_compute34_in[128:65], zll_main_compute34_in[64:1], 3'h2};
  ZLL_Main_compute2  instR10 (zll_main_compute2_inR2[130:67], zll_main_compute2_inR2[66:3], zll_main_compute2_inR2[2:0], zll_main_compute2_outR2);
  assign zll_main_compute2_inR3 = {zll_main_compute34_in[128:65], zll_main_compute34_in[64:1], 3'h3};
  ZLL_Main_compute2  instR11 (zll_main_compute2_inR3[130:67], zll_main_compute2_inR3[66:3], zll_main_compute2_inR3[2:0], zll_main_compute2_outR3);
  assign zll_main_compute2_inR4 = {zll_main_compute34_in[128:65], zll_main_compute34_in[64:1], 3'h4};
  ZLL_Main_compute2  instR12 (zll_main_compute2_inR4[130:67], zll_main_compute2_inR4[66:3], zll_main_compute2_inR4[2:0], zll_main_compute2_outR4);
  assign zll_main_compute2_inR5 = {zll_main_compute34_in[128:65], zll_main_compute34_in[64:1], 3'h5};
  ZLL_Main_compute2  instR13 (zll_main_compute2_inR5[130:67], zll_main_compute2_inR5[66:3], zll_main_compute2_inR5[2:0], zll_main_compute2_outR5);
  assign zll_main_compute2_inR6 = {zll_main_compute34_in[128:65], zll_main_compute34_in[64:1], 3'h6};
  ZLL_Main_compute2  instR14 (zll_main_compute2_inR6[130:67], zll_main_compute2_inR6[66:3], zll_main_compute2_inR6[2:0], zll_main_compute2_outR6);
  assign zll_main_compute2_inR7 = {zll_main_compute34_in[128:65], zll_main_compute34_in[64:1], 3'h7};
  ZLL_Main_compute2  instR15 (zll_main_compute2_inR7[130:67], zll_main_compute2_inR7[66:3], zll_main_compute2_inR7[2:0], zll_main_compute2_outR7);
  assign resize_inR11 = {zll_main_compute2_out, zll_main_compute2_outR1, zll_main_compute2_outR2, zll_main_compute2_outR3, zll_main_compute2_outR4, zll_main_compute2_outR5, zll_main_compute2_outR6, zll_main_compute2_outR7};
  assign resize_inR12 = zll_main_compute34_in[131:129];
  assign binop_inR12 = {128'(resize_inR12[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR13 = {binop_inR12[255:128] * binop_inR12[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR13 = binop_inR13[255:128] % binop_inR13[127:0];
  assign resize_inR14 = resize_inR13[2:0];
  assign binop_inR14 = {128'(resize_inR14[2:0]), 128'h00000000000000000000000000000001};
  assign binop_inR15 = {binop_inR14[255:128] + binop_inR14[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR15 = binop_inR15[255:128] % binop_inR15[127:0];
  assign resize_inR16 = resize_inR15[2:0];
  assign binop_inR16 = {128'h00000000000000000000000000000008, 128'(resize_inR16[2:0])};
  assign binop_inR17 = {binop_inR16[255:128] - binop_inR16[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR18 = {binop_inR17[255:128] - binop_inR17[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR19 = {128'(resize_inR11[63:0]), binop_inR18[255:128] * binop_inR18[127:0]};
  assign resize_inR17 = binop_inR19[255:128] >> binop_inR19[127:0];
  assign res = (zll_main_compute34_in[0] == 1'h1) ? resize_inR17[7:0] : resize_inR10[7:0];
endmodule

module ZLL_Main_compute41 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [127:0] resize_inR1;
  logic [0:0] msbit_in;
  logic [0:0] rewire_prelude_not_in;
  logic [0:0] rewire_prelude_not_out;
  logic [2:0] resize_inR2;
  logic [127:0] resize_inR3;
  logic [0:0] msbit_inR1;
  logic [0:0] rewire_prelude_not_inR1;
  logic [0:0] rewire_prelude_not_outR1;
  logic [131:0] zll_main_compute40_in;
  logic [130:0] zll_main_compute39_in;
  logic [7:0] zll_main_compute39_out;
  logic [130:0] zll_main_compute39_inR1;
  logic [7:0] zll_main_compute39_outR1;
  logic [130:0] zll_main_compute39_inR2;
  logic [7:0] zll_main_compute39_outR2;
  logic [130:0] zll_main_compute39_inR3;
  logic [7:0] zll_main_compute39_outR3;
  logic [130:0] zll_main_compute39_inR4;
  logic [7:0] zll_main_compute39_outR4;
  logic [130:0] zll_main_compute39_inR5;
  logic [7:0] zll_main_compute39_outR5;
  logic [130:0] zll_main_compute39_inR6;
  logic [7:0] zll_main_compute39_outR6;
  logic [130:0] zll_main_compute39_inR7;
  logic [7:0] zll_main_compute39_outR7;
  logic [63:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR8;
  logic [2:0] resize_inR9;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR10;
  logic [2:0] resize_inR11;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR12;
  logic [131:0] zll_main_compute30_in;
  logic [130:0] zll_main_compute29_in;
  logic [7:0] zll_main_compute29_out;
  logic [130:0] zll_main_compute29_inR1;
  logic [7:0] zll_main_compute29_outR1;
  logic [130:0] zll_main_compute29_inR2;
  logic [7:0] zll_main_compute29_outR2;
  logic [130:0] zll_main_compute29_inR3;
  logic [7:0] zll_main_compute29_outR3;
  logic [130:0] zll_main_compute29_inR4;
  logic [7:0] zll_main_compute29_outR4;
  logic [130:0] zll_main_compute29_inR5;
  logic [7:0] zll_main_compute29_outR5;
  logic [130:0] zll_main_compute29_inR6;
  logic [7:0] zll_main_compute29_outR6;
  logic [130:0] zll_main_compute29_inR7;
  logic [7:0] zll_main_compute29_outR7;
  logic [63:0] resize_inR13;
  logic [2:0] resize_inR14;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR15;
  logic [2:0] resize_inR16;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [127:0] resize_inR17;
  logic [2:0] resize_inR18;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [255:0] binop_inR16;
  logic [255:0] binop_inR17;
  logic [127:0] resize_inR19;
  assign resize_in = arg2;
  assign resize_inR1 = 128'(resize_in[2:0]);
  assign msbit_in = resize_inR1[0];
  assign rewire_prelude_not_in = msbit_in[0];
  ReWire_Prelude_not  inst (rewire_prelude_not_in[0], rewire_prelude_not_out);
  assign resize_inR2 = arg2;
  assign resize_inR3 = 128'(resize_inR2[2:0]);
  assign msbit_inR1 = resize_inR3[0];
  assign rewire_prelude_not_inR1 = msbit_inR1[0];
  ReWire_Prelude_not  instR1 (rewire_prelude_not_inR1[0], rewire_prelude_not_outR1);
  assign zll_main_compute40_in = {arg0, arg1, arg2, rewire_prelude_not_outR1};
  assign zll_main_compute39_in = {zll_main_compute40_in[131:68], zll_main_compute40_in[67:4], 3'h0};
  ZLL_Main_compute39  instR2 (zll_main_compute39_in[130:67], zll_main_compute39_in[66:3], zll_main_compute39_in[2:0], zll_main_compute39_out);
  assign zll_main_compute39_inR1 = {zll_main_compute40_in[131:68], zll_main_compute40_in[67:4], 3'h1};
  ZLL_Main_compute39  instR3 (zll_main_compute39_inR1[130:67], zll_main_compute39_inR1[66:3], zll_main_compute39_inR1[2:0], zll_main_compute39_outR1);
  assign zll_main_compute39_inR2 = {zll_main_compute40_in[131:68], zll_main_compute40_in[67:4], 3'h2};
  ZLL_Main_compute39  instR4 (zll_main_compute39_inR2[130:67], zll_main_compute39_inR2[66:3], zll_main_compute39_inR2[2:0], zll_main_compute39_outR2);
  assign zll_main_compute39_inR3 = {zll_main_compute40_in[131:68], zll_main_compute40_in[67:4], 3'h3};
  ZLL_Main_compute39  instR5 (zll_main_compute39_inR3[130:67], zll_main_compute39_inR3[66:3], zll_main_compute39_inR3[2:0], zll_main_compute39_outR3);
  assign zll_main_compute39_inR4 = {zll_main_compute40_in[131:68], zll_main_compute40_in[67:4], 3'h4};
  ZLL_Main_compute39  instR6 (zll_main_compute39_inR4[130:67], zll_main_compute39_inR4[66:3], zll_main_compute39_inR4[2:0], zll_main_compute39_outR4);
  assign zll_main_compute39_inR5 = {zll_main_compute40_in[131:68], zll_main_compute40_in[67:4], 3'h5};
  ZLL_Main_compute39  instR7 (zll_main_compute39_inR5[130:67], zll_main_compute39_inR5[66:3], zll_main_compute39_inR5[2:0], zll_main_compute39_outR5);
  assign zll_main_compute39_inR6 = {zll_main_compute40_in[131:68], zll_main_compute40_in[67:4], 3'h6};
  ZLL_Main_compute39  instR8 (zll_main_compute39_inR6[130:67], zll_main_compute39_inR6[66:3], zll_main_compute39_inR6[2:0], zll_main_compute39_outR6);
  assign zll_main_compute39_inR7 = {zll_main_compute40_in[131:68], zll_main_compute40_in[67:4], 3'h7};
  ZLL_Main_compute39  instR9 (zll_main_compute39_inR7[130:67], zll_main_compute39_inR7[66:3], zll_main_compute39_inR7[2:0], zll_main_compute39_outR7);
  assign resize_inR4 = {zll_main_compute39_out, zll_main_compute39_outR1, zll_main_compute39_outR2, zll_main_compute39_outR3, zll_main_compute39_outR4, zll_main_compute39_outR5, zll_main_compute39_outR6, zll_main_compute39_outR7};
  assign resize_inR5 = zll_main_compute40_in[3:1];
  assign binop_in = {128'(resize_inR5[2:0]), 128'h00000000000000000000000000000001};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR6 = binop_inR1[255:128] % binop_inR1[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR2 = {128'h00000000000000000000000000000003, 128'(resize_inR7[2:0])};
  assign binop_inR3 = {binop_inR2[255:128] + binop_inR2[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR8 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR9 = resize_inR8[2:0];
  assign binop_inR4 = {128'(resize_inR9[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR5 = {binop_inR4[255:128] / binop_inR4[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR10 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR11 = resize_inR10[2:0];
  assign binop_inR6 = {128'h00000000000000000000000000000008, 128'(resize_inR11[2:0])};
  assign binop_inR7 = {binop_inR6[255:128] - binop_inR6[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR8 = {binop_inR7[255:128] - binop_inR7[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR9 = {128'(resize_inR4[63:0]), binop_inR8[255:128] * binop_inR8[127:0]};
  assign resize_inR12 = binop_inR9[255:128] >> binop_inR9[127:0];
  assign zll_main_compute30_in = {arg0, arg1, arg2, rewire_prelude_not_out};
  assign zll_main_compute29_in = {zll_main_compute30_in[131:68], zll_main_compute30_in[67:4], 3'h0};
  ZLL_Main_compute29  instR10 (zll_main_compute29_in[130:67], zll_main_compute29_in[66:3], zll_main_compute29_in[2:0], zll_main_compute29_out);
  assign zll_main_compute29_inR1 = {zll_main_compute30_in[131:68], zll_main_compute30_in[67:4], 3'h1};
  ZLL_Main_compute29  instR11 (zll_main_compute29_inR1[130:67], zll_main_compute29_inR1[66:3], zll_main_compute29_inR1[2:0], zll_main_compute29_outR1);
  assign zll_main_compute29_inR2 = {zll_main_compute30_in[131:68], zll_main_compute30_in[67:4], 3'h2};
  ZLL_Main_compute29  instR12 (zll_main_compute29_inR2[130:67], zll_main_compute29_inR2[66:3], zll_main_compute29_inR2[2:0], zll_main_compute29_outR2);
  assign zll_main_compute29_inR3 = {zll_main_compute30_in[131:68], zll_main_compute30_in[67:4], 3'h3};
  ZLL_Main_compute29  instR13 (zll_main_compute29_inR3[130:67], zll_main_compute29_inR3[66:3], zll_main_compute29_inR3[2:0], zll_main_compute29_outR3);
  assign zll_main_compute29_inR4 = {zll_main_compute30_in[131:68], zll_main_compute30_in[67:4], 3'h4};
  ZLL_Main_compute29  instR14 (zll_main_compute29_inR4[130:67], zll_main_compute29_inR4[66:3], zll_main_compute29_inR4[2:0], zll_main_compute29_outR4);
  assign zll_main_compute29_inR5 = {zll_main_compute30_in[131:68], zll_main_compute30_in[67:4], 3'h5};
  ZLL_Main_compute29  instR15 (zll_main_compute29_inR5[130:67], zll_main_compute29_inR5[66:3], zll_main_compute29_inR5[2:0], zll_main_compute29_outR5);
  assign zll_main_compute29_inR6 = {zll_main_compute30_in[131:68], zll_main_compute30_in[67:4], 3'h6};
  ZLL_Main_compute29  instR16 (zll_main_compute29_inR6[130:67], zll_main_compute29_inR6[66:3], zll_main_compute29_inR6[2:0], zll_main_compute29_outR6);
  assign zll_main_compute29_inR7 = {zll_main_compute30_in[131:68], zll_main_compute30_in[67:4], 3'h7};
  ZLL_Main_compute29  instR17 (zll_main_compute29_inR7[130:67], zll_main_compute29_inR7[66:3], zll_main_compute29_inR7[2:0], zll_main_compute29_outR7);
  assign resize_inR13 = {zll_main_compute29_out, zll_main_compute29_outR1, zll_main_compute29_outR2, zll_main_compute29_outR3, zll_main_compute29_outR4, zll_main_compute29_outR5, zll_main_compute29_outR6, zll_main_compute29_outR7};
  assign resize_inR14 = zll_main_compute30_in[3:1];
  assign binop_inR10 = {128'h00000000000000000000000000000003, 128'(resize_inR14[2:0])};
  assign binop_inR11 = {binop_inR10[255:128] + binop_inR10[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR15 = binop_inR11[255:128] % binop_inR11[127:0];
  assign resize_inR16 = resize_inR15[2:0];
  assign binop_inR12 = {128'(resize_inR16[2:0]), 128'h00000000000000000000000000000002};
  assign binop_inR13 = {binop_inR12[255:128] / binop_inR12[127:0], 128'h00000000000000000000000000000008};
  assign resize_inR17 = binop_inR13[255:128] % binop_inR13[127:0];
  assign resize_inR18 = resize_inR17[2:0];
  assign binop_inR14 = {128'h00000000000000000000000000000008, 128'(resize_inR18[2:0])};
  assign binop_inR15 = {binop_inR14[255:128] - binop_inR14[127:0], 128'h00000000000000000000000000000001};
  assign binop_inR16 = {binop_inR15[255:128] - binop_inR15[127:0], 128'h00000000000000000000000000000008};
  assign binop_inR17 = {128'(resize_inR13[63:0]), binop_inR16[255:128] * binop_inR16[127:0]};
  assign resize_inR19 = binop_inR17[255:128] >> binop_inR17[127:0];
  assign res = (zll_main_compute30_in[0] == 1'h1) ? resize_inR19[7:0] : resize_inR12[7:0];
endmodule

module ReWire_Prelude_not (input logic [0:0] arg0,
  output logic [0:0] res);
  logic [0:0] lit_in;
  assign lit_in = arg0;
  assign res = (lit_in[0] == 1'h1) ? 1'h0 : 1'h1;
endmodule