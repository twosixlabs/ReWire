module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [9:0] __in0,
  output logic [15:0] __out0);
  logic [39:0] rewire_monad_iterst_in;
  logic [69:0] zll_rewire_monad_iterst4_in;
  logic [69:0] zll_rewire_monad_iterst26_in;
  logic [39:0] main_loop1_in;
  logic [29:0] id_in;
  logic [24:0] main_inputtomystate_in;
  logic [24:0] zll_main_inputtomystate23_in;
  logic [13:0] zll_main_inputtomystate18_in;
  logic [24:0] zll_main_inputtomystate6_in;
  logic [24:0] zll_main_inputtomystate12_in;
  logic [12:0] zll_main_inputtomystate24_in;
  logic [24:0] zll_main_inputtomystate7_in;
  logic [22:0] zll_main_inputtomystate5_in;
  logic [22:0] zll_main_inputtomystate14_in;
  logic [24:0] zll_main_inputtomystate26_in;
  logic [18:0] zll_main_inputtomystate27_in;
  logic [13:0] zll_main_inputtomystate19_in;
  logic [44:0] main_incrpipeline_in;
  logic [44:0] zll_main_incrpipeline1_in;
  logic [29:0] id_inR1;
  logic [29:0] resize_in;
  logic [255:0] binop_in;
  logic [127:0] resize_inR1;
  logic [44:0] zll_main_loop3_in;
  logic [14:0] main_mystatetooutput_in;
  logic [14:0] zll_main_mystatetooutput1_in;
  logic [8:0] zll_main_mystatetooutput5_in;
  logic [14:0] zll_main_mystatetooutput3_in;
  logic [12:0] zll_main_mystatetooutput_in;
  logic [14:0] zll_main_mystatetooutput4_in;
  logic [8:0] zll_main_mystatetooutput2_in;
  logic [75:0] zll_rewire_monad_iterst10_in;
  logic [75:0] zll_rewire_monad_iterst32_in;
  logic [77:0] zll_rewire_monad_iterst20_in;
  logic [77:0] zll_rewire_monad_iterst35_in;
  logic [75:0] zll_rewire_monad_iterst14_in;
  logic [75:0] zll_rewire_monad_iterst29_in;
  logic [75:0] zll_rewire_monad_iterst38_in;
  logic [75:0] zll_rewire_monad_iterst25_in;
  logic [29:0] zll_rewire_monad_iterst41_in;
  logic [93:0] zll_rewire_monad_iterst30_in;
  logic [93:0] zll_rewire_monad_iterst24_in;
  logic [45:0] zll_rewire_monad_iterst37_in;
  logic [0:0] __continue;
  logic [30:0] __padding;
  logic [29:0] __st0;
  logic [29:0] __st0_next;
  assign rewire_monad_iterst_in = {__in0, __st0};
  assign zll_rewire_monad_iterst4_in = {rewire_monad_iterst_in[39:30], rewire_monad_iterst_in[29:0], rewire_monad_iterst_in[29:0]};
  assign zll_rewire_monad_iterst26_in = {zll_rewire_monad_iterst4_in[69:60], zll_rewire_monad_iterst4_in[59:0]};
  assign main_loop1_in = {zll_rewire_monad_iterst26_in[69:60], zll_rewire_monad_iterst26_in[59:30]};
  assign id_in = main_loop1_in[29:0];
  assign main_inputtomystate_in = {main_loop1_in[39:30], id_in[29:15]};
  assign zll_main_inputtomystate23_in = {main_inputtomystate_in[24:15], main_inputtomystate_in[14:0]};
  assign zll_main_inputtomystate18_in = {zll_main_inputtomystate23_in[13:9], zll_main_inputtomystate23_in[8:0]};
  assign zll_main_inputtomystate6_in = {main_inputtomystate_in[24:15], main_inputtomystate_in[14:0]};
  assign zll_main_inputtomystate12_in = {main_inputtomystate_in[24:15], main_inputtomystate_in[14:0]};
  assign zll_main_inputtomystate24_in = {zll_main_inputtomystate12_in[12:9], zll_main_inputtomystate12_in[8:0]};
  assign zll_main_inputtomystate7_in = {main_inputtomystate_in[24:15], main_inputtomystate_in[14:0]};
  assign zll_main_inputtomystate5_in = {zll_main_inputtomystate7_in[22:15], zll_main_inputtomystate7_in[14], zll_main_inputtomystate7_in[13:9], zll_main_inputtomystate7_in[8:0]};
  assign zll_main_inputtomystate14_in = {zll_main_inputtomystate5_in[13:9], zll_main_inputtomystate5_in[22:15], zll_main_inputtomystate5_in[14], zll_main_inputtomystate5_in[8:0]};
  assign zll_main_inputtomystate26_in = {main_inputtomystate_in[24:15], main_inputtomystate_in[14:0]};
  assign zll_main_inputtomystate27_in = {zll_main_inputtomystate26_in[18:15], zll_main_inputtomystate26_in[14], zll_main_inputtomystate26_in[13:9], zll_main_inputtomystate26_in[8:0]};
  assign zll_main_inputtomystate19_in = {zll_main_inputtomystate27_in[18:15], zll_main_inputtomystate27_in[14], zll_main_inputtomystate27_in[8:0]};
  assign main_incrpipeline_in = {(zll_main_inputtomystate26_in[24:23] == 2'h0) ? {zll_main_inputtomystate19_in[9], 1'h1, zll_main_inputtomystate19_in[13:10], 5'h00, zll_main_inputtomystate19_in[13:10]} : ((zll_main_inputtomystate7_in[24:23] == 2'h1) ? {zll_main_inputtomystate14_in[9], zll_main_inputtomystate14_in[22:18], 1'h1, zll_main_inputtomystate14_in[17:10]} : (((zll_main_inputtomystate12_in[24:23] == 2'h2) && ((zll_main_inputtomystate12_in[15] == 1'h1) && (zll_main_inputtomystate12_in[13] == 1'h1))) ? {11'h400, zll_main_inputtomystate24_in[12:9]} : (((zll_main_inputtomystate6_in[24:23] == 2'h2) && ((zll_main_inputtomystate6_in[15] == 1'h1) && (zll_main_inputtomystate6_in[13] == 1'h0))) ? {6'h20, zll_main_inputtomystate6_in[8:0]} : {6'h00, zll_main_inputtomystate18_in[8:0]}))), main_loop1_in[29:0]};
  assign zll_main_incrpipeline1_in = main_incrpipeline_in[44:0];
  assign id_inR1 = zll_main_incrpipeline1_in[29:0];
  assign resize_in = zll_main_incrpipeline1_in[29:0];
  assign binop_in = {128'(resize_in[29:0]), {8'h80{1'h0}}};
  assign resize_inR1 = binop_in[255:128] >> binop_in[127:0];
  assign zll_main_loop3_in = {zll_main_incrpipeline1_in[44:30], id_inR1[29:15], resize_inR1[14:0]};
  assign main_mystatetooutput_in = zll_main_loop3_in[14:0];
  assign zll_main_mystatetooutput1_in = main_mystatetooutput_in[14:0];
  assign zll_main_mystatetooutput5_in = zll_main_mystatetooutput1_in[8:0];
  assign zll_main_mystatetooutput3_in = main_mystatetooutput_in[14:0];
  assign zll_main_mystatetooutput_in = {zll_main_mystatetooutput3_in[13:9], zll_main_mystatetooutput3_in[7:0]};
  assign zll_main_mystatetooutput4_in = main_mystatetooutput_in[14:0];
  assign zll_main_mystatetooutput2_in = {zll_main_mystatetooutput4_in[13:9], zll_main_mystatetooutput4_in[3:0]};
  assign zll_rewire_monad_iterst10_in = {{((zll_main_mystatetooutput4_in[14] == 1'h1) && (zll_main_mystatetooutput4_in[8] == 1'h0)) ? {2'h3, zll_main_mystatetooutput2_in[8:4], 5'h00, zll_main_mystatetooutput2_in[3:0]} : (((zll_main_mystatetooutput3_in[14] == 1'h1) && (zll_main_mystatetooutput3_in[8] == 1'h1)) ? {2'h1, zll_main_mystatetooutput_in[12:8], 1'h1, zll_main_mystatetooutput_in[7:0]} : {7'h00, zll_main_mystatetooutput5_in[8:0]}), zll_main_loop3_in[44:15]}, zll_rewire_monad_iterst26_in[29:0]};
  assign zll_rewire_monad_iterst32_in = zll_rewire_monad_iterst10_in[75:0];
  assign zll_rewire_monad_iterst20_in = {2'h0, zll_rewire_monad_iterst32_in[75:30], zll_rewire_monad_iterst32_in[29:0]};
  assign zll_rewire_monad_iterst35_in = zll_rewire_monad_iterst20_in[77:0];
  assign zll_rewire_monad_iterst14_in = {zll_rewire_monad_iterst35_in[75:30], zll_rewire_monad_iterst35_in[29:0]};
  assign zll_rewire_monad_iterst29_in = {zll_rewire_monad_iterst14_in[29:0], zll_rewire_monad_iterst14_in[75:30]};
  assign zll_rewire_monad_iterst38_in = {zll_rewire_monad_iterst29_in[45:30], zll_rewire_monad_iterst29_in[75:46], zll_rewire_monad_iterst29_in[29:0]};
  assign zll_rewire_monad_iterst25_in = {zll_rewire_monad_iterst38_in[75:60], zll_rewire_monad_iterst38_in[29:0], zll_rewire_monad_iterst38_in[59:30]};
  assign zll_rewire_monad_iterst41_in = zll_rewire_monad_iterst25_in[59:30];
  assign zll_rewire_monad_iterst30_in = {zll_rewire_monad_iterst25_in[75:60], {{2'h1, {6'h2e{1'h0}}}, zll_rewire_monad_iterst41_in[29:0]}};
  assign zll_rewire_monad_iterst24_in = {zll_rewire_monad_iterst30_in[93:78], zll_rewire_monad_iterst30_in[77:0]};
  assign zll_rewire_monad_iterst37_in = {zll_rewire_monad_iterst24_in[93:78], zll_rewire_monad_iterst24_in[29:0]};
  assign {__continue, __padding, __out0, __st0_next} = {{1'h1, {5'h1f{1'h0}}}, zll_rewire_monad_iterst37_in[45:30], zll_rewire_monad_iterst37_in[29:0]};
  initial __st0 <= 30'h00000000;
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      __st0 <= 30'h00000000;
    end else begin
      __st0 <= __st0_next;
    end
  end
endmodule