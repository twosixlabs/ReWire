module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [16:0] __in0,
  output logic [14:0] __out0);
  logic [90:0] gzdLLzicase17861;
  logic [143:0] callRes;
  logic [90:0] gzdLLzicase17864;
  logic [143:0] callResR1;
  logic [90:0] gzdLLzicase17867;
  logic [143:0] callResR2;
  logic [90:0] gzdLLzicase17870;
  logic [143:0] callResR3;
  logic [90:0] gzdLLzicase17873;
  logic [143:0] callResR4;
  logic [90:0] gzdLLzicase17876;
  logic [143:0] callResR5;
  logic [90:0] gzdLLzicase17879;
  logic [143:0] callResR6;
  logic [90:0] gzdLLzicase17882;
  logic [143:0] callResR7;
  logic [90:0] gzdLLzicase17885;
  logic [143:0] callResR8;
  logic [0:0] __continue;
  logic [53:0] __padding;
  logic [3:0] __resumption_tag;
  logic [69:0] __st0;
  logic [3:0] __resumption_tag_next;
  logic [69:0] __st0_next;
  assign gzdLLzicase17861 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase17861  zdLLzicase17861 (gzdLLzicase17861[86:17], gzdLLzicase17861[16:0], callRes);
  assign gzdLLzicase17864 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase17864  zdLLzicase17864 (gzdLLzicase17864[86:17], gzdLLzicase17864[16:0], callResR1);
  assign gzdLLzicase17867 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase17867  zdLLzicase17867 (gzdLLzicase17867[86:17], gzdLLzicase17867[16:0], callResR2);
  assign gzdLLzicase17870 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase17870  zdLLzicase17870 (gzdLLzicase17870[86:17], gzdLLzicase17870[16:0], callResR3);
  assign gzdLLzicase17873 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase17873  zdLLzicase17873 (gzdLLzicase17873[86:17], gzdLLzicase17873[16:0], callResR4);
  assign gzdLLzicase17876 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase17876  zdLLzicase17876 (gzdLLzicase17876[86:17], gzdLLzicase17876[16:0], callResR5);
  assign gzdLLzicase17879 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase17879  zdLLzicase17879 (gzdLLzicase17879[86:17], gzdLLzicase17879[16:0], callResR6);
  assign gzdLLzicase17882 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase17882  zdLLzicase17882 (gzdLLzicase17882[86:17], gzdLLzicase17882[16:0], callResR7);
  assign gzdLLzicase17885 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase17885  zdLLzicase17885 (gzdLLzicase17885[86:17], gzdLLzicase17885[16:0], callResR8);
  assign {__continue, __padding, __out0, __resumption_tag_next, __st0_next} = (gzdLLzicase17885[90:87] == 4'h0) ? callResR8 : ((gzdLLzicase17882[90:87] == 4'h1) ? callResR7 : ((gzdLLzicase17879[90:87] == 4'h2) ? callResR6 : ((gzdLLzicase17876[90:87] == 4'h3) ? callResR5 : ((gzdLLzicase17873[90:87] == 4'h4) ? callResR4 : ((gzdLLzicase17870[90:87] == 4'h5) ? callResR3 : ((gzdLLzicase17867[90:87] == 4'h6) ? callResR2 : ((gzdLLzicase17864[90:87] == 4'h7) ? callResR1 : callRes)))))));
  initial {__resumption_tag, __st0} <= {1'h1, {7'h49{1'h0}}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      {__resumption_tag, __st0} <= {1'h1, {7'h49{1'h0}}};
    end else begin
      {__resumption_tag, __st0} <= {__resumption_tag_next, __st0_next};
    end
  end
endmodule

module zdLLzicase14914 (input logic [7:0] arg0,
  input logic [7:0] arg1,
  input logic [7:0] arg2,
  input logic [7:0] arg3,
  input logic [5:0] arg4,
  input logic [16:0] arg5,
  input logic [14:0] arg6,
  input logic [5:0] arg7,
  output logic [69:0] res);
  assign res = {arg0, arg1, arg2, arg3, arg7, arg5, arg6};
endmodule

module zdLLzicase14928 (input logic [7:0] arg0,
  input logic [7:0] arg1,
  input logic [7:0] arg2,
  input logic [7:0] arg3,
  input logic [5:0] arg4,
  input logic [16:0] arg5,
  input logic [14:0] arg6,
  input logic [14:0] arg7,
  output logic [69:0] res);
  assign res = {arg0, arg1, arg2, arg3, arg4, arg5, arg7};
endmodule

module zdLLzicase14938 (input logic [0:0] arg0,
  input logic [5:0] arg1,
  input logic [7:0] arg2,
  input logic [5:0] arg3,
  output logic [14:0] res);
  assign res = {arg0, arg3, arg2};
endmodule

module zdLLzicase14964 (input logic [0:0] arg0,
  input logic [5:0] arg1,
  input logic [7:0] arg2,
  output logic [14:0] res);
  assign res = {1'h0, arg1, arg2};
endmodule

module zdLLzicase14973 (input logic [7:0] arg0,
  input logic [7:0] arg1,
  input logic [7:0] arg2,
  input logic [7:0] arg3,
  input logic [5:0] arg4,
  input logic [16:0] arg5,
  input logic [14:0] arg6,
  input logic [16:0] arg7,
  output logic [69:0] res);
  assign res = {arg0, arg1, arg2, arg3, arg4, arg7, arg6};
endmodule

module zdLLzicase15143 (input logic [7:0] arg0,
  input logic [7:0] arg1,
  input logic [7:0] arg2,
  input logic [7:0] arg3,
  input logic [5:0] arg4,
  input logic [16:0] arg5,
  input logic [14:0] arg6,
  input logic [7:0] arg7,
  output logic [69:0] res);
  assign res = {arg7, arg1, arg2, arg3, arg4, arg5, arg6};
endmodule

module zdLLzicase17861 (input logic [69:0] arg0,
  input logic [16:0] arg1,
  output logic [143:0] res);
  logic [86:0] gzdLLzilambda16190;
  logic [86:0] gzdLLzilambda16107;
  logic [139:0] gzdLLzilambda19317;
  logic [139:0] gzdLLzicase18021;
  logic [143:0] callRes;
  logic [160:0] gzdLLzilambda19312;
  logic [160:0] gzdLLzicase19309;
  logic [156:0] gzdLLzilambda16105;
  logic [86:0] gzdLLzicase14973;
  logic [69:0] callResR1;
  logic [69:0] gzdLLzicase17968;
  logic [143:0] callResR2;
  logic [143:0] gzdLLzilambda19452;
  logic [143:0] gzdLLzicase19450;
  logic [69:0] gzdLLzilambda16188;
  logic [139:0] gzdLLzilambda19447;
  logic [139:0] gzdLLzicase18021R1;
  logic [143:0] callResR3;
  logic [143:0] gzdLLzilambda19442;
  logic [143:0] gzdLLzicase19440;
  logic [139:0] gzdLLzilambda16186;
  logic [69:0] gMainzipc;
  logic [5:0] callResR4;
  logic [143:0] gzdLLzilambda19437;
  logic [143:0] gzdLLzicase19435;
  logic [75:0] gzdLLzilambda16184;
  logic [75:0] gzdLLzilambda16134;
  logic [139:0] gzdLLzilambda19353;
  logic [139:0] gzdLLzicase18021R2;
  logic [143:0] callResR5;
  logic [149:0] gzdLLzilambda19348;
  logic [149:0] gzdLLzicase19345;
  logic [145:0] gzdLLzilambda16132;
  logic [69:0] gMainzioutputs;
  logic [14:0] callResR6;
  logic [149:0] gzdLLzilambda19341;
  logic [149:0] gzdLLzicase19338;
  logic [90:0] gzdLLzilambda16129;
  logic [20:0] gzdLLzicase14938;
  logic [14:0] callResR7;
  logic [84:0] gzdLLzilambda16121;
  logic [139:0] gzdLLzilambda19334;
  logic [139:0] gzdLLzicase18021R3;
  logic [143:0] callResR8;
  logic [158:0] gzdLLzilambda19329;
  logic [158:0] gzdLLzicase19326;
  logic [154:0] gzdLLzilambda16119;
  logic [84:0] gzdLLzicase14928;
  logic [69:0] callResR9;
  logic [69:0] gzdLLzicase17968R1;
  logic [143:0] callResR10;
  logic [143:0] gzdLLzilambda19432;
  logic [143:0] gzdLLzicase19430;
  logic [69:0] gzdLLzilambda16182;
  logic [139:0] gzdLLzilambda19427;
  logic [139:0] gzdLLzicase18021R4;
  logic [143:0] callResR11;
  logic [143:0] gzdLLzilambda19422;
  logic [143:0] gzdLLzicase19420;
  logic [139:0] gzdLLzilambda16180;
  logic [69:0] gMainzioutputsR1;
  logic [14:0] callResR12;
  logic [143:0] gzdLLzilambda19417;
  logic [143:0] gzdLLzicase19415;
  logic [84:0] gzdLLzilambda16178;
  logic [14:0] gzdLLzicase14964;
  logic [14:0] callResR13;
  logic [84:0] gzdLLzilambda16148;
  logic [139:0] gzdLLzilambda19370;
  logic [139:0] gzdLLzicase18021R5;
  logic [143:0] callResR14;
  logic [158:0] gzdLLzilambda19365;
  logic [158:0] gzdLLzicase19362;
  logic [154:0] gzdLLzilambda16146;
  logic [84:0] gzdLLzicase14928R1;
  logic [69:0] callResR15;
  logic [69:0] gzdLLzicase17968R2;
  logic [143:0] callResR16;
  logic [143:0] gzdLLzilambda19412;
  logic [143:0] gzdLLzicase19410;
  logic [69:0] gzdLLzilambda16176;
  logic [139:0] gzdLLzilambda19407;
  logic [139:0] gzdLLzicase18021R6;
  logic [143:0] callResR17;
  logic [143:0] gzdLLzilambda19402;
  logic [143:0] gzdLLzicase19400;
  logic [139:0] gzdLLzilambda16174;
  logic [69:0] gMainzioutputsR2;
  logic [14:0] callResR18;
  logic [143:0] gzdLLzilambda19397;
  logic [143:0] gzdLLzicase19395;
  logic [84:0] gzdLLzilambda16172;
  assign gzdLLzilambda16190 = {arg1, arg0};
  assign gzdLLzilambda16107 = {gzdLLzilambda16190[86:70], gzdLLzilambda16190[69:0]};
  assign gzdLLzilambda19317 = {gzdLLzilambda16107[69:0], gzdLLzilambda16107[69:0]};
  assign gzdLLzicase18021 = gzdLLzilambda19317[139:0];
  zdLLzicase18021  zdLLzicase18021 (gzdLLzicase18021[139:70], gzdLLzicase18021[69:0], callRes);
  assign gzdLLzilambda19312 = {gzdLLzilambda16107[86:70], callRes};
  assign gzdLLzicase19309 = {gzdLLzilambda19312[143:0], gzdLLzilambda19312[160:144]};
  assign gzdLLzilambda16105 = {gzdLLzicase19309[16:0], gzdLLzicase19309[156:87], gzdLLzicase19309[86:17]};
  assign gzdLLzicase14973 = {gzdLLzilambda16105[139:70], gzdLLzilambda16105[156:140]};
  zdLLzicase14973  zdLLzicase14973 (gzdLLzicase14973[86:79], gzdLLzicase14973[78:71], gzdLLzicase14973[70:63], gzdLLzicase14973[62:55], gzdLLzicase14973[54:49], gzdLLzicase14973[48:32], gzdLLzicase14973[31:17], gzdLLzicase14973[16:0], callResR1);
  assign gzdLLzicase17968 = callResR1;
  zdLLzicase17968  zdLLzicase17968 (gzdLLzicase17968[69:0], callResR2);
  assign gzdLLzilambda19452 = callResR2;
  assign gzdLLzicase19450 = gzdLLzilambda19452[143:0];
  assign gzdLLzilambda16188 = gzdLLzicase19450[69:0];
  assign gzdLLzilambda19447 = {gzdLLzilambda16188[69:0], gzdLLzilambda16188[69:0]};
  assign gzdLLzicase18021R1 = gzdLLzilambda19447[139:0];
  zdLLzicase18021  zdLLzicase18021R1 (gzdLLzicase18021R1[139:70], gzdLLzicase18021R1[69:0], callResR3);
  assign gzdLLzilambda19442 = callResR3;
  assign gzdLLzicase19440 = gzdLLzilambda19442[143:0];
  assign gzdLLzilambda16186 = {gzdLLzicase19440[139:70], gzdLLzicase19440[69:0]};
  assign gMainzipc = gzdLLzilambda16186[139:70];
  Mainzipc  Mainzipc (gMainzipc[69:0], callResR4);
  assign gzdLLzilambda19437 = {{7'h44{1'h0}}, callResR4, gzdLLzilambda16186[69:0]};
  assign gzdLLzicase19435 = gzdLLzilambda19437[143:0];
  assign gzdLLzilambda16184 = {gzdLLzicase19435[75:70], gzdLLzicase19435[69:0]};
  assign gzdLLzilambda16134 = {gzdLLzilambda16184[75:70], gzdLLzilambda16184[69:0]};
  assign gzdLLzilambda19353 = {gzdLLzilambda16134[69:0], gzdLLzilambda16134[69:0]};
  assign gzdLLzicase18021R2 = gzdLLzilambda19353[139:0];
  zdLLzicase18021  zdLLzicase18021R2 (gzdLLzicase18021R2[139:70], gzdLLzicase18021R2[69:0], callResR5);
  assign gzdLLzilambda19348 = {gzdLLzilambda16134[75:70], callResR5};
  assign gzdLLzicase19345 = {gzdLLzilambda19348[143:0], gzdLLzilambda19348[149:144]};
  assign gzdLLzilambda16132 = {gzdLLzicase19345[5:0], gzdLLzicase19345[145:76], gzdLLzicase19345[75:6]};
  assign gMainzioutputs = gzdLLzilambda16132[139:70];
  Mainzioutputs  Mainzioutputs (gMainzioutputs[69:0], callResR6);
  assign gzdLLzilambda19341 = {gzdLLzilambda16132[145:140], {4'h5, {6'h37{1'h0}}}, callResR6, gzdLLzilambda16132[69:0]};
  assign gzdLLzicase19338 = {gzdLLzilambda19341[143:0], gzdLLzilambda19341[149:144]};
  assign gzdLLzilambda16129 = {gzdLLzicase19338[5:0], gzdLLzicase19338[90:76], gzdLLzicase19338[75:6]};
  assign gzdLLzicase14938 = {gzdLLzilambda16129[84:70], gzdLLzilambda16129[90:85]};
  zdLLzicase14938  zdLLzicase14938 (gzdLLzicase14938[20], gzdLLzicase14938[19:14], gzdLLzicase14938[13:6], gzdLLzicase14938[5:0], callResR7);
  assign gzdLLzilambda16121 = {callResR7, gzdLLzilambda16129[69:0]};
  assign gzdLLzilambda19334 = {gzdLLzilambda16121[69:0], gzdLLzilambda16121[69:0]};
  assign gzdLLzicase18021R3 = gzdLLzilambda19334[139:0];
  zdLLzicase18021  zdLLzicase18021R3 (gzdLLzicase18021R3[139:70], gzdLLzicase18021R3[69:0], callResR8);
  assign gzdLLzilambda19329 = {gzdLLzilambda16121[84:70], callResR8};
  assign gzdLLzicase19326 = {gzdLLzilambda19329[143:0], gzdLLzilambda19329[158:144]};
  assign gzdLLzilambda16119 = {gzdLLzicase19326[14:0], gzdLLzicase19326[154:85], gzdLLzicase19326[84:15]};
  assign gzdLLzicase14928 = {gzdLLzilambda16119[139:70], gzdLLzilambda16119[154:140]};
  zdLLzicase14928  zdLLzicase14928 (gzdLLzicase14928[84:77], gzdLLzicase14928[76:69], gzdLLzicase14928[68:61], gzdLLzicase14928[60:53], gzdLLzicase14928[52:47], gzdLLzicase14928[46:30], gzdLLzicase14928[29:15], gzdLLzicase14928[14:0], callResR9);
  assign gzdLLzicase17968R1 = callResR9;
  zdLLzicase17968  zdLLzicase17968R1 (gzdLLzicase17968R1[69:0], callResR10);
  assign gzdLLzilambda19432 = callResR10;
  assign gzdLLzicase19430 = gzdLLzilambda19432[143:0];
  assign gzdLLzilambda16182 = gzdLLzicase19430[69:0];
  assign gzdLLzilambda19427 = {gzdLLzilambda16182[69:0], gzdLLzilambda16182[69:0]};
  assign gzdLLzicase18021R4 = gzdLLzilambda19427[139:0];
  zdLLzicase18021  zdLLzicase18021R4 (gzdLLzicase18021R4[139:70], gzdLLzicase18021R4[69:0], callResR11);
  assign gzdLLzilambda19422 = callResR11;
  assign gzdLLzicase19420 = gzdLLzilambda19422[143:0];
  assign gzdLLzilambda16180 = {gzdLLzicase19420[139:70], gzdLLzicase19420[69:0]};
  assign gMainzioutputsR1 = gzdLLzilambda16180[139:70];
  Mainzioutputs  MainzioutputsR1 (gMainzioutputsR1[69:0], callResR12);
  assign gzdLLzilambda19417 = {{4'h5, {6'h37{1'h0}}}, callResR12, gzdLLzilambda16180[69:0]};
  assign gzdLLzicase19415 = gzdLLzilambda19417[143:0];
  assign gzdLLzilambda16178 = {gzdLLzicase19415[84:70], gzdLLzicase19415[69:0]};
  assign gzdLLzicase14964 = gzdLLzilambda16178[84:70];
  zdLLzicase14964  zdLLzicase14964 (gzdLLzicase14964[14], gzdLLzicase14964[13:8], gzdLLzicase14964[7:0], callResR13);
  assign gzdLLzilambda16148 = {callResR13, gzdLLzilambda16178[69:0]};
  assign gzdLLzilambda19370 = {gzdLLzilambda16148[69:0], gzdLLzilambda16148[69:0]};
  assign gzdLLzicase18021R5 = gzdLLzilambda19370[139:0];
  zdLLzicase18021  zdLLzicase18021R5 (gzdLLzicase18021R5[139:70], gzdLLzicase18021R5[69:0], callResR14);
  assign gzdLLzilambda19365 = {gzdLLzilambda16148[84:70], callResR14};
  assign gzdLLzicase19362 = {gzdLLzilambda19365[143:0], gzdLLzilambda19365[158:144]};
  assign gzdLLzilambda16146 = {gzdLLzicase19362[14:0], gzdLLzicase19362[154:85], gzdLLzicase19362[84:15]};
  assign gzdLLzicase14928R1 = {gzdLLzilambda16146[139:70], gzdLLzilambda16146[154:140]};
  zdLLzicase14928  zdLLzicase14928R1 (gzdLLzicase14928R1[84:77], gzdLLzicase14928R1[76:69], gzdLLzicase14928R1[68:61], gzdLLzicase14928R1[60:53], gzdLLzicase14928R1[52:47], gzdLLzicase14928R1[46:30], gzdLLzicase14928R1[29:15], gzdLLzicase14928R1[14:0], callResR15);
  assign gzdLLzicase17968R2 = callResR15;
  zdLLzicase17968  zdLLzicase17968R2 (gzdLLzicase17968R2[69:0], callResR16);
  assign gzdLLzilambda19412 = callResR16;
  assign gzdLLzicase19410 = gzdLLzilambda19412[143:0];
  assign gzdLLzilambda16176 = gzdLLzicase19410[69:0];
  assign gzdLLzilambda19407 = {gzdLLzilambda16176[69:0], gzdLLzilambda16176[69:0]};
  assign gzdLLzicase18021R6 = gzdLLzilambda19407[139:0];
  zdLLzicase18021  zdLLzicase18021R6 (gzdLLzicase18021R6[139:70], gzdLLzicase18021R6[69:0], callResR17);
  assign gzdLLzilambda19402 = callResR17;
  assign gzdLLzicase19400 = gzdLLzilambda19402[143:0];
  assign gzdLLzilambda16174 = {gzdLLzicase19400[139:70], gzdLLzicase19400[69:0]};
  assign gMainzioutputsR2 = gzdLLzilambda16174[139:70];
  Mainzioutputs  MainzioutputsR2 (gMainzioutputsR2[69:0], callResR18);
  assign gzdLLzilambda19397 = {{4'h5, {6'h37{1'h0}}}, callResR18, gzdLLzilambda16174[69:0]};
  assign gzdLLzicase19395 = gzdLLzilambda19397[143:0];
  assign gzdLLzilambda16172 = {gzdLLzicase19395[84:70], gzdLLzicase19395[69:0]};
  assign res = {{1'h1, {6'h36{1'h0}}}, gzdLLzilambda16172[84:70], 4'h7, gzdLLzilambda16172[69:0]};
endmodule

module zdLLzicase17864 (input logic [69:0] arg0,
  input logic [16:0] arg1,
  output logic [143:0] res);
  logic [86:0] gzdLLzilambda16170;
  logic [86:0] gzdLLzilambda16166;
  logic [139:0] gzdLLzilambda19387;
  logic [139:0] gzdLLzicase18021;
  logic [143:0] callRes;
  logic [160:0] gzdLLzilambda19382;
  logic [160:0] gzdLLzicase19379;
  logic [156:0] gzdLLzilambda16164;
  logic [86:0] gzdLLzicase14973;
  logic [69:0] callResR1;
  logic [69:0] gzdLLzicase17968;
  logic [143:0] callResR2;
  logic [143:0] gzdLLzilambda19392;
  logic [143:0] gzdLLzicase19243;
  logic [143:0] callResR3;
  assign gzdLLzilambda16170 = {arg1, arg0};
  assign gzdLLzilambda16166 = {gzdLLzilambda16170[86:70], gzdLLzilambda16170[69:0]};
  assign gzdLLzilambda19387 = {gzdLLzilambda16166[69:0], gzdLLzilambda16166[69:0]};
  assign gzdLLzicase18021 = gzdLLzilambda19387[139:0];
  zdLLzicase18021  zdLLzicase18021 (gzdLLzicase18021[139:70], gzdLLzicase18021[69:0], callRes);
  assign gzdLLzilambda19382 = {gzdLLzilambda16166[86:70], callRes};
  assign gzdLLzicase19379 = {gzdLLzilambda19382[143:0], gzdLLzilambda19382[160:144]};
  assign gzdLLzilambda16164 = {gzdLLzicase19379[16:0], gzdLLzicase19379[156:87], gzdLLzicase19379[86:17]};
  assign gzdLLzicase14973 = {gzdLLzilambda16164[139:70], gzdLLzilambda16164[156:140]};
  zdLLzicase14973  zdLLzicase14973 (gzdLLzicase14973[86:79], gzdLLzicase14973[78:71], gzdLLzicase14973[70:63], gzdLLzicase14973[62:55], gzdLLzicase14973[54:49], gzdLLzicase14973[48:32], gzdLLzicase14973[31:17], gzdLLzicase14973[16:0], callResR1);
  assign gzdLLzicase17968 = callResR1;
  zdLLzicase17968  zdLLzicase17968 (gzdLLzicase17968[69:0], callResR2);
  assign gzdLLzilambda19392 = callResR2;
  assign gzdLLzicase19243 = gzdLLzilambda19392[143:0];
  zdLLzicase19243  zdLLzicase19243 (gzdLLzicase19243[69:0], callResR3);
  assign res = callResR3;
endmodule

module zdLLzicase17867 (input logic [69:0] arg0,
  input logic [16:0] arg1,
  output logic [143:0] res);
  logic [86:0] gzdLLzilambda15708;
  logic [139:0] gzdLLzilambda19158;
  logic [139:0] gzdLLzicase18021;
  logic [143:0] callRes;
  logic [160:0] gzdLLzilambda19153;
  logic [160:0] gzdLLzicase19150;
  logic [156:0] gzdLLzilambda15706;
  logic [86:0] gzdLLzicase14973;
  logic [69:0] callResR1;
  logic [69:0] gzdLLzicase17968;
  logic [143:0] callResR2;
  assign gzdLLzilambda15708 = {arg1, arg0};
  assign gzdLLzilambda19158 = {gzdLLzilambda15708[69:0], gzdLLzilambda15708[69:0]};
  assign gzdLLzicase18021 = gzdLLzilambda19158[139:0];
  zdLLzicase18021  zdLLzicase18021 (gzdLLzicase18021[139:70], gzdLLzicase18021[69:0], callRes);
  assign gzdLLzilambda19153 = {gzdLLzilambda15708[86:70], callRes};
  assign gzdLLzicase19150 = {gzdLLzilambda19153[143:0], gzdLLzilambda19153[160:144]};
  assign gzdLLzilambda15706 = {gzdLLzicase19150[16:0], gzdLLzicase19150[156:87], gzdLLzicase19150[86:17]};
  assign gzdLLzicase14973 = {gzdLLzilambda15706[139:70], gzdLLzilambda15706[156:140]};
  zdLLzicase14973  zdLLzicase14973 (gzdLLzicase14973[86:79], gzdLLzicase14973[78:71], gzdLLzicase14973[70:63], gzdLLzicase14973[62:55], gzdLLzicase14973[54:49], gzdLLzicase14973[48:32], gzdLLzicase14973[31:17], gzdLLzicase14973[16:0], callResR1);
  assign gzdLLzicase17968 = callResR1;
  zdLLzicase17968  zdLLzicase17968 (gzdLLzicase17968[69:0], callResR2);
  assign res = callResR2;
endmodule

module zdLLzicase17870 (input logic [69:0] arg0,
  input logic [16:0] arg1,
  output logic [143:0] res);
  logic [86:0] gzdLLzilambda15569;
  logic [139:0] gzdLLzilambda18951;
  logic [139:0] gzdLLzicase18021;
  logic [143:0] callRes;
  logic [160:0] gzdLLzilambda18946;
  logic [160:0] gzdLLzicase18943;
  logic [156:0] gzdLLzilambda15567;
  logic [86:0] gzdLLzicase14973;
  logic [69:0] callResR1;
  logic [69:0] gzdLLzicase17968;
  logic [143:0] callResR2;
  assign gzdLLzilambda15569 = {arg1, arg0};
  assign gzdLLzilambda18951 = {gzdLLzilambda15569[69:0], gzdLLzilambda15569[69:0]};
  assign gzdLLzicase18021 = gzdLLzilambda18951[139:0];
  zdLLzicase18021  zdLLzicase18021 (gzdLLzicase18021[139:70], gzdLLzicase18021[69:0], callRes);
  assign gzdLLzilambda18946 = {gzdLLzilambda15569[86:70], callRes};
  assign gzdLLzicase18943 = {gzdLLzilambda18946[143:0], gzdLLzilambda18946[160:144]};
  assign gzdLLzilambda15567 = {gzdLLzicase18943[16:0], gzdLLzicase18943[156:87], gzdLLzicase18943[86:17]};
  assign gzdLLzicase14973 = {gzdLLzilambda15567[139:70], gzdLLzilambda15567[156:140]};
  zdLLzicase14973  zdLLzicase14973 (gzdLLzicase14973[86:79], gzdLLzicase14973[78:71], gzdLLzicase14973[70:63], gzdLLzicase14973[62:55], gzdLLzicase14973[54:49], gzdLLzicase14973[48:32], gzdLLzicase14973[31:17], gzdLLzicase14973[16:0], callResR1);
  assign gzdLLzicase17968 = callResR1;
  zdLLzicase17968  zdLLzicase17968 (gzdLLzicase17968[69:0], callResR2);
  assign res = callResR2;
endmodule

module zdLLzicase17873 (input logic [69:0] arg0,
  input logic [16:0] arg1,
  output logic [143:0] res);
  logic [86:0] gzdLLzilambda15387;
  logic [86:0] gzdLLzilambda15286;
  logic [139:0] gzdLLzilambda18605;
  logic [139:0] gzdLLzicase18021;
  logic [143:0] callRes;
  logic [160:0] gzdLLzilambda18600;
  logic [160:0] gzdLLzicase18597;
  logic [156:0] gzdLLzilambda15284;
  logic [86:0] gzdLLzicase14973;
  logic [69:0] callResR1;
  logic [69:0] gzdLLzicase17968;
  logic [143:0] callResR2;
  logic [143:0] gzdLLzilambda18772;
  logic [143:0] gzdLLzicase18770;
  logic [69:0] gzdLLzilambda15385;
  logic [139:0] gzdLLzilambda18767;
  logic [139:0] gzdLLzicase18021R1;
  logic [143:0] callResR3;
  logic [143:0] gzdLLzilambda18762;
  logic [143:0] gzdLLzicase18760;
  logic [139:0] gzdLLzilambda15383;
  logic [69:0] gMainzipc;
  logic [5:0] callResR4;
  logic [143:0] gzdLLzilambda18757;
  logic [143:0] gzdLLzicase18755;
  logic [75:0] gzdLLzilambda15381;
  logic [11:0] binOp;
  logic [75:0] gzdLLzilambda15300;
  logic [139:0] gzdLLzilambda18622;
  logic [139:0] gzdLLzicase18021R2;
  logic [143:0] callResR5;
  logic [149:0] gzdLLzilambda18617;
  logic [149:0] gzdLLzicase18614;
  logic [145:0] gzdLLzilambda15298;
  logic [75:0] gzdLLzicase14914;
  logic [69:0] callResR6;
  logic [69:0] gzdLLzicase17968R1;
  logic [143:0] callResR7;
  logic [143:0] gzdLLzilambda18752;
  logic [143:0] gzdLLzicase18750;
  logic [69:0] gzdLLzilambda15379;
  logic [139:0] gzdLLzilambda18747;
  logic [139:0] gzdLLzicase18021R3;
  logic [143:0] callResR8;
  logic [143:0] gzdLLzilambda18742;
  logic [143:0] gzdLLzicase18740;
  logic [139:0] gzdLLzilambda15377;
  logic [69:0] gMainzipcR1;
  logic [5:0] callResR9;
  logic [143:0] gzdLLzilambda18737;
  logic [143:0] gzdLLzicase18735;
  logic [75:0] gzdLLzilambda15375;
  logic [75:0] gzdLLzilambda15327;
  logic [139:0] gzdLLzilambda18658;
  logic [139:0] gzdLLzicase18021R4;
  logic [143:0] callResR10;
  logic [149:0] gzdLLzilambda18653;
  logic [149:0] gzdLLzicase18650;
  logic [145:0] gzdLLzilambda15325;
  logic [69:0] gMainzioutputs;
  logic [14:0] callResR11;
  logic [149:0] gzdLLzilambda18646;
  logic [149:0] gzdLLzicase18643;
  logic [90:0] gzdLLzilambda15322;
  logic [20:0] gzdLLzicase14938;
  logic [14:0] callResR12;
  logic [84:0] gzdLLzilambda15314;
  logic [139:0] gzdLLzilambda18639;
  logic [139:0] gzdLLzicase18021R5;
  logic [143:0] callResR13;
  logic [158:0] gzdLLzilambda18634;
  logic [158:0] gzdLLzicase18631;
  logic [154:0] gzdLLzilambda15312;
  logic [84:0] gzdLLzicase14928;
  logic [69:0] callResR14;
  logic [69:0] gzdLLzicase17968R2;
  logic [143:0] callResR15;
  logic [143:0] gzdLLzilambda18732;
  logic [143:0] gzdLLzicase18730;
  logic [69:0] gzdLLzilambda15373;
  logic [139:0] gzdLLzilambda18727;
  logic [139:0] gzdLLzicase18021R6;
  logic [143:0] callResR16;
  logic [143:0] gzdLLzilambda18722;
  logic [143:0] gzdLLzicase18720;
  logic [139:0] gzdLLzilambda15371;
  logic [69:0] gMainzioutputsR1;
  logic [14:0] callResR17;
  logic [143:0] gzdLLzilambda18717;
  logic [143:0] gzdLLzicase18715;
  logic [84:0] gzdLLzilambda15369;
  logic [14:0] gzdLLzicase14964;
  logic [14:0] callResR18;
  logic [84:0] gzdLLzilambda15341;
  logic [139:0] gzdLLzilambda18675;
  logic [139:0] gzdLLzicase18021R7;
  logic [143:0] callResR19;
  logic [158:0] gzdLLzilambda18670;
  logic [158:0] gzdLLzicase18667;
  logic [154:0] gzdLLzilambda15339;
  logic [84:0] gzdLLzicase14928R1;
  logic [69:0] callResR20;
  logic [69:0] gzdLLzicase17968R3;
  logic [143:0] callResR21;
  logic [143:0] gzdLLzilambda18712;
  logic [143:0] gzdLLzicase18710;
  logic [69:0] gzdLLzilambda15367;
  logic [139:0] gzdLLzilambda18707;
  logic [139:0] gzdLLzicase18021R8;
  logic [143:0] callResR22;
  logic [143:0] gzdLLzilambda18702;
  logic [143:0] gzdLLzicase18700;
  logic [139:0] gzdLLzilambda15365;
  logic [69:0] gMainzioutputsR2;
  logic [14:0] callResR23;
  logic [143:0] gzdLLzilambda18697;
  logic [143:0] gzdLLzicase18695;
  logic [84:0] gzdLLzilambda15363;
  assign gzdLLzilambda15387 = {arg1, arg0};
  assign gzdLLzilambda15286 = {gzdLLzilambda15387[86:70], gzdLLzilambda15387[69:0]};
  assign gzdLLzilambda18605 = {gzdLLzilambda15286[69:0], gzdLLzilambda15286[69:0]};
  assign gzdLLzicase18021 = gzdLLzilambda18605[139:0];
  zdLLzicase18021  zdLLzicase18021 (gzdLLzicase18021[139:70], gzdLLzicase18021[69:0], callRes);
  assign gzdLLzilambda18600 = {gzdLLzilambda15286[86:70], callRes};
  assign gzdLLzicase18597 = {gzdLLzilambda18600[143:0], gzdLLzilambda18600[160:144]};
  assign gzdLLzilambda15284 = {gzdLLzicase18597[16:0], gzdLLzicase18597[156:87], gzdLLzicase18597[86:17]};
  assign gzdLLzicase14973 = {gzdLLzilambda15284[139:70], gzdLLzilambda15284[156:140]};
  zdLLzicase14973  zdLLzicase14973 (gzdLLzicase14973[86:79], gzdLLzicase14973[78:71], gzdLLzicase14973[70:63], gzdLLzicase14973[62:55], gzdLLzicase14973[54:49], gzdLLzicase14973[48:32], gzdLLzicase14973[31:17], gzdLLzicase14973[16:0], callResR1);
  assign gzdLLzicase17968 = callResR1;
  zdLLzicase17968  zdLLzicase17968 (gzdLLzicase17968[69:0], callResR2);
  assign gzdLLzilambda18772 = callResR2;
  assign gzdLLzicase18770 = gzdLLzilambda18772[143:0];
  assign gzdLLzilambda15385 = gzdLLzicase18770[69:0];
  assign gzdLLzilambda18767 = {gzdLLzilambda15385[69:0], gzdLLzilambda15385[69:0]};
  assign gzdLLzicase18021R1 = gzdLLzilambda18767[139:0];
  zdLLzicase18021  zdLLzicase18021R1 (gzdLLzicase18021R1[139:70], gzdLLzicase18021R1[69:0], callResR3);
  assign gzdLLzilambda18762 = callResR3;
  assign gzdLLzicase18760 = gzdLLzilambda18762[143:0];
  assign gzdLLzilambda15383 = {gzdLLzicase18760[139:70], gzdLLzicase18760[69:0]};
  assign gMainzipc = gzdLLzilambda15383[139:70];
  Mainzipc  Mainzipc (gMainzipc[69:0], callResR4);
  assign gzdLLzilambda18757 = {{7'h44{1'h0}}, callResR4, gzdLLzilambda15383[69:0]};
  assign gzdLLzicase18755 = gzdLLzilambda18757[143:0];
  assign gzdLLzilambda15381 = {gzdLLzicase18755[75:70], gzdLLzicase18755[69:0]};
  assign binOp = {gzdLLzilambda15381[75:70], 6'h01};
  assign gzdLLzilambda15300 = {binOp[11:6] + binOp[5:0], gzdLLzilambda15381[69:0]};
  assign gzdLLzilambda18622 = {gzdLLzilambda15300[69:0], gzdLLzilambda15300[69:0]};
  assign gzdLLzicase18021R2 = gzdLLzilambda18622[139:0];
  zdLLzicase18021  zdLLzicase18021R2 (gzdLLzicase18021R2[139:70], gzdLLzicase18021R2[69:0], callResR5);
  assign gzdLLzilambda18617 = {gzdLLzilambda15300[75:70], callResR5};
  assign gzdLLzicase18614 = {gzdLLzilambda18617[143:0], gzdLLzilambda18617[149:144]};
  assign gzdLLzilambda15298 = {gzdLLzicase18614[5:0], gzdLLzicase18614[145:76], gzdLLzicase18614[75:6]};
  assign gzdLLzicase14914 = {gzdLLzilambda15298[139:70], gzdLLzilambda15298[145:140]};
  zdLLzicase14914  zdLLzicase14914 (gzdLLzicase14914[75:68], gzdLLzicase14914[67:60], gzdLLzicase14914[59:52], gzdLLzicase14914[51:44], gzdLLzicase14914[43:38], gzdLLzicase14914[37:21], gzdLLzicase14914[20:6], gzdLLzicase14914[5:0], callResR6);
  assign gzdLLzicase17968R1 = callResR6;
  zdLLzicase17968  zdLLzicase17968R1 (gzdLLzicase17968R1[69:0], callResR7);
  assign gzdLLzilambda18752 = callResR7;
  assign gzdLLzicase18750 = gzdLLzilambda18752[143:0];
  assign gzdLLzilambda15379 = gzdLLzicase18750[69:0];
  assign gzdLLzilambda18747 = {gzdLLzilambda15379[69:0], gzdLLzilambda15379[69:0]};
  assign gzdLLzicase18021R3 = gzdLLzilambda18747[139:0];
  zdLLzicase18021  zdLLzicase18021R3 (gzdLLzicase18021R3[139:70], gzdLLzicase18021R3[69:0], callResR8);
  assign gzdLLzilambda18742 = callResR8;
  assign gzdLLzicase18740 = gzdLLzilambda18742[143:0];
  assign gzdLLzilambda15377 = {gzdLLzicase18740[139:70], gzdLLzicase18740[69:0]};
  assign gMainzipcR1 = gzdLLzilambda15377[139:70];
  Mainzipc  MainzipcR1 (gMainzipcR1[69:0], callResR9);
  assign gzdLLzilambda18737 = {{7'h44{1'h0}}, callResR9, gzdLLzilambda15377[69:0]};
  assign gzdLLzicase18735 = gzdLLzilambda18737[143:0];
  assign gzdLLzilambda15375 = {gzdLLzicase18735[75:70], gzdLLzicase18735[69:0]};
  assign gzdLLzilambda15327 = {gzdLLzilambda15375[75:70], gzdLLzilambda15375[69:0]};
  assign gzdLLzilambda18658 = {gzdLLzilambda15327[69:0], gzdLLzilambda15327[69:0]};
  assign gzdLLzicase18021R4 = gzdLLzilambda18658[139:0];
  zdLLzicase18021  zdLLzicase18021R4 (gzdLLzicase18021R4[139:70], gzdLLzicase18021R4[69:0], callResR10);
  assign gzdLLzilambda18653 = {gzdLLzilambda15327[75:70], callResR10};
  assign gzdLLzicase18650 = {gzdLLzilambda18653[143:0], gzdLLzilambda18653[149:144]};
  assign gzdLLzilambda15325 = {gzdLLzicase18650[5:0], gzdLLzicase18650[145:76], gzdLLzicase18650[75:6]};
  assign gMainzioutputs = gzdLLzilambda15325[139:70];
  Mainzioutputs  Mainzioutputs (gMainzioutputs[69:0], callResR11);
  assign gzdLLzilambda18646 = {gzdLLzilambda15325[145:140], {4'h5, {6'h37{1'h0}}}, callResR11, gzdLLzilambda15325[69:0]};
  assign gzdLLzicase18643 = {gzdLLzilambda18646[143:0], gzdLLzilambda18646[149:144]};
  assign gzdLLzilambda15322 = {gzdLLzicase18643[5:0], gzdLLzicase18643[90:76], gzdLLzicase18643[75:6]};
  assign gzdLLzicase14938 = {gzdLLzilambda15322[84:70], gzdLLzilambda15322[90:85]};
  zdLLzicase14938  zdLLzicase14938 (gzdLLzicase14938[20], gzdLLzicase14938[19:14], gzdLLzicase14938[13:6], gzdLLzicase14938[5:0], callResR12);
  assign gzdLLzilambda15314 = {callResR12, gzdLLzilambda15322[69:0]};
  assign gzdLLzilambda18639 = {gzdLLzilambda15314[69:0], gzdLLzilambda15314[69:0]};
  assign gzdLLzicase18021R5 = gzdLLzilambda18639[139:0];
  zdLLzicase18021  zdLLzicase18021R5 (gzdLLzicase18021R5[139:70], gzdLLzicase18021R5[69:0], callResR13);
  assign gzdLLzilambda18634 = {gzdLLzilambda15314[84:70], callResR13};
  assign gzdLLzicase18631 = {gzdLLzilambda18634[143:0], gzdLLzilambda18634[158:144]};
  assign gzdLLzilambda15312 = {gzdLLzicase18631[14:0], gzdLLzicase18631[154:85], gzdLLzicase18631[84:15]};
  assign gzdLLzicase14928 = {gzdLLzilambda15312[139:70], gzdLLzilambda15312[154:140]};
  zdLLzicase14928  zdLLzicase14928 (gzdLLzicase14928[84:77], gzdLLzicase14928[76:69], gzdLLzicase14928[68:61], gzdLLzicase14928[60:53], gzdLLzicase14928[52:47], gzdLLzicase14928[46:30], gzdLLzicase14928[29:15], gzdLLzicase14928[14:0], callResR14);
  assign gzdLLzicase17968R2 = callResR14;
  zdLLzicase17968  zdLLzicase17968R2 (gzdLLzicase17968R2[69:0], callResR15);
  assign gzdLLzilambda18732 = callResR15;
  assign gzdLLzicase18730 = gzdLLzilambda18732[143:0];
  assign gzdLLzilambda15373 = gzdLLzicase18730[69:0];
  assign gzdLLzilambda18727 = {gzdLLzilambda15373[69:0], gzdLLzilambda15373[69:0]};
  assign gzdLLzicase18021R6 = gzdLLzilambda18727[139:0];
  zdLLzicase18021  zdLLzicase18021R6 (gzdLLzicase18021R6[139:70], gzdLLzicase18021R6[69:0], callResR16);
  assign gzdLLzilambda18722 = callResR16;
  assign gzdLLzicase18720 = gzdLLzilambda18722[143:0];
  assign gzdLLzilambda15371 = {gzdLLzicase18720[139:70], gzdLLzicase18720[69:0]};
  assign gMainzioutputsR1 = gzdLLzilambda15371[139:70];
  Mainzioutputs  MainzioutputsR1 (gMainzioutputsR1[69:0], callResR17);
  assign gzdLLzilambda18717 = {{4'h5, {6'h37{1'h0}}}, callResR17, gzdLLzilambda15371[69:0]};
  assign gzdLLzicase18715 = gzdLLzilambda18717[143:0];
  assign gzdLLzilambda15369 = {gzdLLzicase18715[84:70], gzdLLzicase18715[69:0]};
  assign gzdLLzicase14964 = gzdLLzilambda15369[84:70];
  zdLLzicase14964  zdLLzicase14964 (gzdLLzicase14964[14], gzdLLzicase14964[13:8], gzdLLzicase14964[7:0], callResR18);
  assign gzdLLzilambda15341 = {callResR18, gzdLLzilambda15369[69:0]};
  assign gzdLLzilambda18675 = {gzdLLzilambda15341[69:0], gzdLLzilambda15341[69:0]};
  assign gzdLLzicase18021R7 = gzdLLzilambda18675[139:0];
  zdLLzicase18021  zdLLzicase18021R7 (gzdLLzicase18021R7[139:70], gzdLLzicase18021R7[69:0], callResR19);
  assign gzdLLzilambda18670 = {gzdLLzilambda15341[84:70], callResR19};
  assign gzdLLzicase18667 = {gzdLLzilambda18670[143:0], gzdLLzilambda18670[158:144]};
  assign gzdLLzilambda15339 = {gzdLLzicase18667[14:0], gzdLLzicase18667[154:85], gzdLLzicase18667[84:15]};
  assign gzdLLzicase14928R1 = {gzdLLzilambda15339[139:70], gzdLLzilambda15339[154:140]};
  zdLLzicase14928  zdLLzicase14928R1 (gzdLLzicase14928R1[84:77], gzdLLzicase14928R1[76:69], gzdLLzicase14928R1[68:61], gzdLLzicase14928R1[60:53], gzdLLzicase14928R1[52:47], gzdLLzicase14928R1[46:30], gzdLLzicase14928R1[29:15], gzdLLzicase14928R1[14:0], callResR20);
  assign gzdLLzicase17968R3 = callResR20;
  zdLLzicase17968  zdLLzicase17968R3 (gzdLLzicase17968R3[69:0], callResR21);
  assign gzdLLzilambda18712 = callResR21;
  assign gzdLLzicase18710 = gzdLLzilambda18712[143:0];
  assign gzdLLzilambda15367 = gzdLLzicase18710[69:0];
  assign gzdLLzilambda18707 = {gzdLLzilambda15367[69:0], gzdLLzilambda15367[69:0]};
  assign gzdLLzicase18021R8 = gzdLLzilambda18707[139:0];
  zdLLzicase18021  zdLLzicase18021R8 (gzdLLzicase18021R8[139:70], gzdLLzicase18021R8[69:0], callResR22);
  assign gzdLLzilambda18702 = callResR22;
  assign gzdLLzicase18700 = gzdLLzilambda18702[143:0];
  assign gzdLLzilambda15365 = {gzdLLzicase18700[139:70], gzdLLzicase18700[69:0]};
  assign gMainzioutputsR2 = gzdLLzilambda15365[139:70];
  Mainzioutputs  MainzioutputsR2 (gMainzioutputsR2[69:0], callResR23);
  assign gzdLLzilambda18697 = {{4'h5, {6'h37{1'h0}}}, callResR23, gzdLLzilambda15365[69:0]};
  assign gzdLLzicase18695 = gzdLLzilambda18697[143:0];
  assign gzdLLzilambda15363 = {gzdLLzicase18695[84:70], gzdLLzicase18695[69:0]};
  assign res = {{1'h1, {6'h36{1'h0}}}, gzdLLzilambda15363[84:70], 4'h3, gzdLLzilambda15363[69:0]};
endmodule

module zdLLzicase17876 (input logic [69:0] arg0,
  input logic [16:0] arg1,
  output logic [143:0] res);
  logic [86:0] gzdLLzilambda15359;
  logic [139:0] gzdLLzilambda18692;
  logic [139:0] gzdLLzicase18021;
  logic [143:0] callRes;
  logic [160:0] gzdLLzilambda18687;
  logic [160:0] gzdLLzicase18684;
  logic [156:0] gzdLLzilambda15357;
  logic [86:0] gzdLLzicase14973;
  logic [69:0] callResR1;
  logic [69:0] gzdLLzicase17968;
  logic [143:0] callResR2;
  assign gzdLLzilambda15359 = {arg1, arg0};
  assign gzdLLzilambda18692 = {gzdLLzilambda15359[69:0], gzdLLzilambda15359[69:0]};
  assign gzdLLzicase18021 = gzdLLzilambda18692[139:0];
  zdLLzicase18021  zdLLzicase18021 (gzdLLzicase18021[139:70], gzdLLzicase18021[69:0], callRes);
  assign gzdLLzilambda18687 = {gzdLLzilambda15359[86:70], callRes};
  assign gzdLLzicase18684 = {gzdLLzilambda18687[143:0], gzdLLzilambda18687[160:144]};
  assign gzdLLzilambda15357 = {gzdLLzicase18684[16:0], gzdLLzicase18684[156:87], gzdLLzicase18684[86:17]};
  assign gzdLLzicase14973 = {gzdLLzilambda15357[139:70], gzdLLzilambda15357[156:140]};
  zdLLzicase14973  zdLLzicase14973 (gzdLLzicase14973[86:79], gzdLLzicase14973[78:71], gzdLLzicase14973[70:63], gzdLLzicase14973[62:55], gzdLLzicase14973[54:49], gzdLLzicase14973[48:32], gzdLLzicase14973[31:17], gzdLLzicase14973[16:0], callResR1);
  assign gzdLLzicase17968 = callResR1;
  zdLLzicase17968  zdLLzicase17968 (gzdLLzicase17968[69:0], callResR2);
  assign res = callResR2;
endmodule

module zdLLzicase17879 (input logic [69:0] arg0,
  input logic [16:0] arg1,
  output logic [143:0] res);
  logic [86:0] gzdLLzilambda15184;
  logic [86:0] gzdLLzilambda15061;
  logic [139:0] gzdLLzilambda18255;
  logic [139:0] gzdLLzicase18021;
  logic [143:0] callRes;
  logic [160:0] gzdLLzilambda18250;
  logic [160:0] gzdLLzicase18247;
  logic [156:0] gzdLLzilambda15059;
  logic [86:0] gzdLLzicase14973;
  logic [69:0] callResR1;
  logic [69:0] gzdLLzicase17968;
  logic [143:0] callResR2;
  logic [143:0] gzdLLzilambda18459;
  logic [143:0] gzdLLzicase18457;
  logic [69:0] gzdLLzilambda15182;
  logic [139:0] gzdLLzilambda18454;
  logic [139:0] gzdLLzicase18021R1;
  logic [143:0] callResR3;
  logic [143:0] gzdLLzilambda18449;
  logic [143:0] gzdLLzicase18447;
  logic [139:0] gzdLLzilambda15180;
  logic [69:0] gMainzipc;
  logic [5:0] callResR4;
  logic [143:0] gzdLLzilambda18444;
  logic [143:0] gzdLLzicase18442;
  logic [75:0] gzdLLzilambda15178;
  logic [11:0] binOp;
  logic [75:0] gzdLLzilambda15075;
  logic [139:0] gzdLLzilambda18272;
  logic [139:0] gzdLLzicase18021R2;
  logic [143:0] callResR5;
  logic [149:0] gzdLLzilambda18267;
  logic [149:0] gzdLLzicase18264;
  logic [145:0] gzdLLzilambda15073;
  logic [75:0] gzdLLzicase14914;
  logic [69:0] callResR6;
  logic [69:0] gzdLLzicase17968R1;
  logic [143:0] callResR7;
  logic [143:0] gzdLLzilambda18439;
  logic [143:0] gzdLLzicase18437;
  logic [69:0] gzdLLzilambda15176;
  logic [139:0] gzdLLzilambda18434;
  logic [139:0] gzdLLzicase18021R3;
  logic [143:0] callResR8;
  logic [143:0] gzdLLzilambda18429;
  logic [143:0] gzdLLzicase18427;
  logic [139:0] gzdLLzilambda15174;
  logic [69:0] gMainzipcR1;
  logic [5:0] callResR9;
  logic [143:0] gzdLLzilambda18424;
  logic [143:0] gzdLLzicase18422;
  logic [75:0] gzdLLzilambda15172;
  logic [75:0] gzdLLzilambda15102;
  logic [139:0] gzdLLzilambda18308;
  logic [139:0] gzdLLzicase18021R4;
  logic [143:0] callResR10;
  logic [149:0] gzdLLzilambda18303;
  logic [149:0] gzdLLzicase18300;
  logic [145:0] gzdLLzilambda15100;
  logic [69:0] gMainzioutputs;
  logic [14:0] callResR11;
  logic [149:0] gzdLLzilambda18296;
  logic [149:0] gzdLLzicase18293;
  logic [90:0] gzdLLzilambda15097;
  logic [20:0] gzdLLzicase14938;
  logic [14:0] callResR12;
  logic [84:0] gzdLLzilambda15089;
  logic [139:0] gzdLLzilambda18289;
  logic [139:0] gzdLLzicase18021R5;
  logic [143:0] callResR13;
  logic [158:0] gzdLLzilambda18284;
  logic [158:0] gzdLLzicase18281;
  logic [154:0] gzdLLzilambda15087;
  logic [84:0] gzdLLzicase14928;
  logic [69:0] callResR14;
  logic [69:0] gzdLLzicase17968R2;
  logic [143:0] callResR15;
  logic [143:0] gzdLLzilambda18419;
  logic [143:0] gzdLLzicase18417;
  logic [69:0] gzdLLzilambda15170;
  logic [139:0] gzdLLzilambda18414;
  logic [139:0] gzdLLzicase18021R6;
  logic [143:0] callResR16;
  logic [143:0] gzdLLzilambda18409;
  logic [143:0] gzdLLzicase18407;
  logic [139:0] gzdLLzilambda15168;
  logic [69:0] gMainzioutputsR1;
  logic [14:0] callResR17;
  logic [143:0] gzdLLzilambda18404;
  logic [143:0] gzdLLzicase18402;
  logic [84:0] gzdLLzilambda15166;
  logic [14:0] gzdLLzicase14964;
  logic [14:0] callResR18;
  logic [84:0] gzdLLzilambda15116;
  logic [139:0] gzdLLzilambda18325;
  logic [139:0] gzdLLzicase18021R7;
  logic [143:0] callResR19;
  logic [158:0] gzdLLzilambda18320;
  logic [158:0] gzdLLzicase18317;
  logic [154:0] gzdLLzilambda15114;
  logic [84:0] gzdLLzicase14928R1;
  logic [69:0] callResR20;
  logic [69:0] gzdLLzicase17968R3;
  logic [143:0] callResR21;
  logic [143:0] gzdLLzilambda18399;
  logic [143:0] gzdLLzicase18397;
  logic [69:0] gzdLLzilambda15164;
  logic [139:0] gzdLLzilambda18394;
  logic [139:0] gzdLLzicase18021R8;
  logic [143:0] callResR22;
  logic [143:0] gzdLLzilambda18389;
  logic [143:0] gzdLLzicase18387;
  logic [139:0] gzdLLzilambda15162;
  logic [69:0] gMainzioutputsR2;
  logic [14:0] callResR23;
  logic [143:0] gzdLLzilambda18384;
  logic [143:0] gzdLLzicase18382;
  logic [84:0] gzdLLzilambda15160;
  assign gzdLLzilambda15184 = {arg1, arg0};
  assign gzdLLzilambda15061 = {gzdLLzilambda15184[86:70], gzdLLzilambda15184[69:0]};
  assign gzdLLzilambda18255 = {gzdLLzilambda15061[69:0], gzdLLzilambda15061[69:0]};
  assign gzdLLzicase18021 = gzdLLzilambda18255[139:0];
  zdLLzicase18021  zdLLzicase18021 (gzdLLzicase18021[139:70], gzdLLzicase18021[69:0], callRes);
  assign gzdLLzilambda18250 = {gzdLLzilambda15061[86:70], callRes};
  assign gzdLLzicase18247 = {gzdLLzilambda18250[143:0], gzdLLzilambda18250[160:144]};
  assign gzdLLzilambda15059 = {gzdLLzicase18247[16:0], gzdLLzicase18247[156:87], gzdLLzicase18247[86:17]};
  assign gzdLLzicase14973 = {gzdLLzilambda15059[139:70], gzdLLzilambda15059[156:140]};
  zdLLzicase14973  zdLLzicase14973 (gzdLLzicase14973[86:79], gzdLLzicase14973[78:71], gzdLLzicase14973[70:63], gzdLLzicase14973[62:55], gzdLLzicase14973[54:49], gzdLLzicase14973[48:32], gzdLLzicase14973[31:17], gzdLLzicase14973[16:0], callResR1);
  assign gzdLLzicase17968 = callResR1;
  zdLLzicase17968  zdLLzicase17968 (gzdLLzicase17968[69:0], callResR2);
  assign gzdLLzilambda18459 = callResR2;
  assign gzdLLzicase18457 = gzdLLzilambda18459[143:0];
  assign gzdLLzilambda15182 = gzdLLzicase18457[69:0];
  assign gzdLLzilambda18454 = {gzdLLzilambda15182[69:0], gzdLLzilambda15182[69:0]};
  assign gzdLLzicase18021R1 = gzdLLzilambda18454[139:0];
  zdLLzicase18021  zdLLzicase18021R1 (gzdLLzicase18021R1[139:70], gzdLLzicase18021R1[69:0], callResR3);
  assign gzdLLzilambda18449 = callResR3;
  assign gzdLLzicase18447 = gzdLLzilambda18449[143:0];
  assign gzdLLzilambda15180 = {gzdLLzicase18447[139:70], gzdLLzicase18447[69:0]};
  assign gMainzipc = gzdLLzilambda15180[139:70];
  Mainzipc  Mainzipc (gMainzipc[69:0], callResR4);
  assign gzdLLzilambda18444 = {{7'h44{1'h0}}, callResR4, gzdLLzilambda15180[69:0]};
  assign gzdLLzicase18442 = gzdLLzilambda18444[143:0];
  assign gzdLLzilambda15178 = {gzdLLzicase18442[75:70], gzdLLzicase18442[69:0]};
  assign binOp = {gzdLLzilambda15178[75:70], 6'h01};
  assign gzdLLzilambda15075 = {binOp[11:6] + binOp[5:0], gzdLLzilambda15178[69:0]};
  assign gzdLLzilambda18272 = {gzdLLzilambda15075[69:0], gzdLLzilambda15075[69:0]};
  assign gzdLLzicase18021R2 = gzdLLzilambda18272[139:0];
  zdLLzicase18021  zdLLzicase18021R2 (gzdLLzicase18021R2[139:70], gzdLLzicase18021R2[69:0], callResR5);
  assign gzdLLzilambda18267 = {gzdLLzilambda15075[75:70], callResR5};
  assign gzdLLzicase18264 = {gzdLLzilambda18267[143:0], gzdLLzilambda18267[149:144]};
  assign gzdLLzilambda15073 = {gzdLLzicase18264[5:0], gzdLLzicase18264[145:76], gzdLLzicase18264[75:6]};
  assign gzdLLzicase14914 = {gzdLLzilambda15073[139:70], gzdLLzilambda15073[145:140]};
  zdLLzicase14914  zdLLzicase14914 (gzdLLzicase14914[75:68], gzdLLzicase14914[67:60], gzdLLzicase14914[59:52], gzdLLzicase14914[51:44], gzdLLzicase14914[43:38], gzdLLzicase14914[37:21], gzdLLzicase14914[20:6], gzdLLzicase14914[5:0], callResR6);
  assign gzdLLzicase17968R1 = callResR6;
  zdLLzicase17968  zdLLzicase17968R1 (gzdLLzicase17968R1[69:0], callResR7);
  assign gzdLLzilambda18439 = callResR7;
  assign gzdLLzicase18437 = gzdLLzilambda18439[143:0];
  assign gzdLLzilambda15176 = gzdLLzicase18437[69:0];
  assign gzdLLzilambda18434 = {gzdLLzilambda15176[69:0], gzdLLzilambda15176[69:0]};
  assign gzdLLzicase18021R3 = gzdLLzilambda18434[139:0];
  zdLLzicase18021  zdLLzicase18021R3 (gzdLLzicase18021R3[139:70], gzdLLzicase18021R3[69:0], callResR8);
  assign gzdLLzilambda18429 = callResR8;
  assign gzdLLzicase18427 = gzdLLzilambda18429[143:0];
  assign gzdLLzilambda15174 = {gzdLLzicase18427[139:70], gzdLLzicase18427[69:0]};
  assign gMainzipcR1 = gzdLLzilambda15174[139:70];
  Mainzipc  MainzipcR1 (gMainzipcR1[69:0], callResR9);
  assign gzdLLzilambda18424 = {{7'h44{1'h0}}, callResR9, gzdLLzilambda15174[69:0]};
  assign gzdLLzicase18422 = gzdLLzilambda18424[143:0];
  assign gzdLLzilambda15172 = {gzdLLzicase18422[75:70], gzdLLzicase18422[69:0]};
  assign gzdLLzilambda15102 = {gzdLLzilambda15172[75:70], gzdLLzilambda15172[69:0]};
  assign gzdLLzilambda18308 = {gzdLLzilambda15102[69:0], gzdLLzilambda15102[69:0]};
  assign gzdLLzicase18021R4 = gzdLLzilambda18308[139:0];
  zdLLzicase18021  zdLLzicase18021R4 (gzdLLzicase18021R4[139:70], gzdLLzicase18021R4[69:0], callResR10);
  assign gzdLLzilambda18303 = {gzdLLzilambda15102[75:70], callResR10};
  assign gzdLLzicase18300 = {gzdLLzilambda18303[143:0], gzdLLzilambda18303[149:144]};
  assign gzdLLzilambda15100 = {gzdLLzicase18300[5:0], gzdLLzicase18300[145:76], gzdLLzicase18300[75:6]};
  assign gMainzioutputs = gzdLLzilambda15100[139:70];
  Mainzioutputs  Mainzioutputs (gMainzioutputs[69:0], callResR11);
  assign gzdLLzilambda18296 = {gzdLLzilambda15100[145:140], {4'h5, {6'h37{1'h0}}}, callResR11, gzdLLzilambda15100[69:0]};
  assign gzdLLzicase18293 = {gzdLLzilambda18296[143:0], gzdLLzilambda18296[149:144]};
  assign gzdLLzilambda15097 = {gzdLLzicase18293[5:0], gzdLLzicase18293[90:76], gzdLLzicase18293[75:6]};
  assign gzdLLzicase14938 = {gzdLLzilambda15097[84:70], gzdLLzilambda15097[90:85]};
  zdLLzicase14938  zdLLzicase14938 (gzdLLzicase14938[20], gzdLLzicase14938[19:14], gzdLLzicase14938[13:6], gzdLLzicase14938[5:0], callResR12);
  assign gzdLLzilambda15089 = {callResR12, gzdLLzilambda15097[69:0]};
  assign gzdLLzilambda18289 = {gzdLLzilambda15089[69:0], gzdLLzilambda15089[69:0]};
  assign gzdLLzicase18021R5 = gzdLLzilambda18289[139:0];
  zdLLzicase18021  zdLLzicase18021R5 (gzdLLzicase18021R5[139:70], gzdLLzicase18021R5[69:0], callResR13);
  assign gzdLLzilambda18284 = {gzdLLzilambda15089[84:70], callResR13};
  assign gzdLLzicase18281 = {gzdLLzilambda18284[143:0], gzdLLzilambda18284[158:144]};
  assign gzdLLzilambda15087 = {gzdLLzicase18281[14:0], gzdLLzicase18281[154:85], gzdLLzicase18281[84:15]};
  assign gzdLLzicase14928 = {gzdLLzilambda15087[139:70], gzdLLzilambda15087[154:140]};
  zdLLzicase14928  zdLLzicase14928 (gzdLLzicase14928[84:77], gzdLLzicase14928[76:69], gzdLLzicase14928[68:61], gzdLLzicase14928[60:53], gzdLLzicase14928[52:47], gzdLLzicase14928[46:30], gzdLLzicase14928[29:15], gzdLLzicase14928[14:0], callResR14);
  assign gzdLLzicase17968R2 = callResR14;
  zdLLzicase17968  zdLLzicase17968R2 (gzdLLzicase17968R2[69:0], callResR15);
  assign gzdLLzilambda18419 = callResR15;
  assign gzdLLzicase18417 = gzdLLzilambda18419[143:0];
  assign gzdLLzilambda15170 = gzdLLzicase18417[69:0];
  assign gzdLLzilambda18414 = {gzdLLzilambda15170[69:0], gzdLLzilambda15170[69:0]};
  assign gzdLLzicase18021R6 = gzdLLzilambda18414[139:0];
  zdLLzicase18021  zdLLzicase18021R6 (gzdLLzicase18021R6[139:70], gzdLLzicase18021R6[69:0], callResR16);
  assign gzdLLzilambda18409 = callResR16;
  assign gzdLLzicase18407 = gzdLLzilambda18409[143:0];
  assign gzdLLzilambda15168 = {gzdLLzicase18407[139:70], gzdLLzicase18407[69:0]};
  assign gMainzioutputsR1 = gzdLLzilambda15168[139:70];
  Mainzioutputs  MainzioutputsR1 (gMainzioutputsR1[69:0], callResR17);
  assign gzdLLzilambda18404 = {{4'h5, {6'h37{1'h0}}}, callResR17, gzdLLzilambda15168[69:0]};
  assign gzdLLzicase18402 = gzdLLzilambda18404[143:0];
  assign gzdLLzilambda15166 = {gzdLLzicase18402[84:70], gzdLLzicase18402[69:0]};
  assign gzdLLzicase14964 = gzdLLzilambda15166[84:70];
  zdLLzicase14964  zdLLzicase14964 (gzdLLzicase14964[14], gzdLLzicase14964[13:8], gzdLLzicase14964[7:0], callResR18);
  assign gzdLLzilambda15116 = {callResR18, gzdLLzilambda15166[69:0]};
  assign gzdLLzilambda18325 = {gzdLLzilambda15116[69:0], gzdLLzilambda15116[69:0]};
  assign gzdLLzicase18021R7 = gzdLLzilambda18325[139:0];
  zdLLzicase18021  zdLLzicase18021R7 (gzdLLzicase18021R7[139:70], gzdLLzicase18021R7[69:0], callResR19);
  assign gzdLLzilambda18320 = {gzdLLzilambda15116[84:70], callResR19};
  assign gzdLLzicase18317 = {gzdLLzilambda18320[143:0], gzdLLzilambda18320[158:144]};
  assign gzdLLzilambda15114 = {gzdLLzicase18317[14:0], gzdLLzicase18317[154:85], gzdLLzicase18317[84:15]};
  assign gzdLLzicase14928R1 = {gzdLLzilambda15114[139:70], gzdLLzilambda15114[154:140]};
  zdLLzicase14928  zdLLzicase14928R1 (gzdLLzicase14928R1[84:77], gzdLLzicase14928R1[76:69], gzdLLzicase14928R1[68:61], gzdLLzicase14928R1[60:53], gzdLLzicase14928R1[52:47], gzdLLzicase14928R1[46:30], gzdLLzicase14928R1[29:15], gzdLLzicase14928R1[14:0], callResR20);
  assign gzdLLzicase17968R3 = callResR20;
  zdLLzicase17968  zdLLzicase17968R3 (gzdLLzicase17968R3[69:0], callResR21);
  assign gzdLLzilambda18399 = callResR21;
  assign gzdLLzicase18397 = gzdLLzilambda18399[143:0];
  assign gzdLLzilambda15164 = gzdLLzicase18397[69:0];
  assign gzdLLzilambda18394 = {gzdLLzilambda15164[69:0], gzdLLzilambda15164[69:0]};
  assign gzdLLzicase18021R8 = gzdLLzilambda18394[139:0];
  zdLLzicase18021  zdLLzicase18021R8 (gzdLLzicase18021R8[139:70], gzdLLzicase18021R8[69:0], callResR22);
  assign gzdLLzilambda18389 = callResR22;
  assign gzdLLzicase18387 = gzdLLzilambda18389[143:0];
  assign gzdLLzilambda15162 = {gzdLLzicase18387[139:70], gzdLLzicase18387[69:0]};
  assign gMainzioutputsR2 = gzdLLzilambda15162[139:70];
  Mainzioutputs  MainzioutputsR2 (gMainzioutputsR2[69:0], callResR23);
  assign gzdLLzilambda18384 = {{4'h5, {6'h37{1'h0}}}, callResR23, gzdLLzilambda15162[69:0]};
  assign gzdLLzicase18382 = gzdLLzilambda18384[143:0];
  assign gzdLLzilambda15160 = {gzdLLzicase18382[84:70], gzdLLzicase18382[69:0]};
  assign res = {{1'h1, {6'h36{1'h0}}}, gzdLLzilambda15160[84:70], 4'h1, gzdLLzilambda15160[69:0]};
endmodule

module zdLLzicase17882 (input logic [69:0] arg0,
  input logic [16:0] arg1,
  output logic [143:0] res);
  logic [86:0] gzdLLzilambda15158;
  logic [86:0] gzdLLzilambda15134;
  logic [139:0] gzdLLzilambda18342;
  logic [139:0] gzdLLzicase18021;
  logic [143:0] callRes;
  logic [160:0] gzdLLzilambda18337;
  logic [160:0] gzdLLzicase18334;
  logic [156:0] gzdLLzilambda15132;
  logic [86:0] gzdLLzicase14973;
  logic [69:0] callResR1;
  logic [69:0] gzdLLzicase17968;
  logic [143:0] callResR2;
  logic [143:0] gzdLLzilambda18379;
  logic [143:0] gzdLLzicase18377;
  logic [69:0] gzdLLzilambda15156;
  logic [139:0] gzdLLzilambda18374;
  logic [139:0] gzdLLzicase18021R1;
  logic [143:0] callResR3;
  logic [143:0] gzdLLzilambda18369;
  logic [143:0] gzdLLzicase18367;
  logic [139:0] gzdLLzilambda15154;
  logic [69:0] gMainziinputs;
  logic [16:0] callResR4;
  logic [143:0] gzdLLzilambda18364;
  logic [143:0] gzdLLzicase18362;
  logic [86:0] gzdLLzilambda15152;
  logic [16:0] gMainzidataIn;
  logic [16:0] gzdLLzicase14627;
  logic [143:0] gzdLLzilambda18359;
  logic [143:0] gzdLLzicase18357;
  logic [77:0] gzdLLzilambda15148;
  logic [147:0] gzdLLzilambda18354;
  logic [147:0] gzdLLzicase18351;
  logic [147:0] gzdLLzilambda15146;
  logic [77:0] gzdLLzicase15143;
  logic [69:0] callResR5;
  logic [69:0] gzdLLzicase17968R1;
  logic [143:0] callResR6;
  assign gzdLLzilambda15158 = {arg1, arg0};
  assign gzdLLzilambda15134 = {gzdLLzilambda15158[86:70], gzdLLzilambda15158[69:0]};
  assign gzdLLzilambda18342 = {gzdLLzilambda15134[69:0], gzdLLzilambda15134[69:0]};
  assign gzdLLzicase18021 = gzdLLzilambda18342[139:0];
  zdLLzicase18021  zdLLzicase18021 (gzdLLzicase18021[139:70], gzdLLzicase18021[69:0], callRes);
  assign gzdLLzilambda18337 = {gzdLLzilambda15134[86:70], callRes};
  assign gzdLLzicase18334 = {gzdLLzilambda18337[143:0], gzdLLzilambda18337[160:144]};
  assign gzdLLzilambda15132 = {gzdLLzicase18334[16:0], gzdLLzicase18334[156:87], gzdLLzicase18334[86:17]};
  assign gzdLLzicase14973 = {gzdLLzilambda15132[139:70], gzdLLzilambda15132[156:140]};
  zdLLzicase14973  zdLLzicase14973 (gzdLLzicase14973[86:79], gzdLLzicase14973[78:71], gzdLLzicase14973[70:63], gzdLLzicase14973[62:55], gzdLLzicase14973[54:49], gzdLLzicase14973[48:32], gzdLLzicase14973[31:17], gzdLLzicase14973[16:0], callResR1);
  assign gzdLLzicase17968 = callResR1;
  zdLLzicase17968  zdLLzicase17968 (gzdLLzicase17968[69:0], callResR2);
  assign gzdLLzilambda18379 = callResR2;
  assign gzdLLzicase18377 = gzdLLzilambda18379[143:0];
  assign gzdLLzilambda15156 = gzdLLzicase18377[69:0];
  assign gzdLLzilambda18374 = {gzdLLzilambda15156[69:0], gzdLLzilambda15156[69:0]};
  assign gzdLLzicase18021R1 = gzdLLzilambda18374[139:0];
  zdLLzicase18021  zdLLzicase18021R1 (gzdLLzicase18021R1[139:70], gzdLLzicase18021R1[69:0], callResR3);
  assign gzdLLzilambda18369 = callResR3;
  assign gzdLLzicase18367 = gzdLLzilambda18369[143:0];
  assign gzdLLzilambda15154 = {gzdLLzicase18367[139:70], gzdLLzicase18367[69:0]};
  assign gMainziinputs = gzdLLzilambda15154[139:70];
  Mainziinputs  Mainziinputs (gMainziinputs[69:0], callResR4);
  assign gzdLLzilambda18364 = {{4'h3, {6'h35{1'h0}}}, callResR4, gzdLLzilambda15154[69:0]};
  assign gzdLLzicase18362 = gzdLLzilambda18364[143:0];
  assign gzdLLzilambda15152 = {gzdLLzicase18362[86:70], gzdLLzicase18362[69:0]};
  assign gMainzidataIn = gzdLLzilambda15152[86:70];
  assign gzdLLzicase14627 = gMainzidataIn[16:0];
  assign gzdLLzilambda18359 = {{4'h1, {6'h3e{1'h0}}}, gzdLLzicase14627[7:0], gzdLLzilambda15152[69:0]};
  assign gzdLLzicase18357 = gzdLLzilambda18359[143:0];
  assign gzdLLzilambda15148 = {gzdLLzicase18357[77:70], gzdLLzicase18357[69:0]};
  assign gzdLLzilambda18354 = {gzdLLzilambda15148[77:70], gzdLLzilambda15148[69:0], gzdLLzilambda15148[69:0]};
  assign gzdLLzicase18351 = {gzdLLzilambda18354[139:0], gzdLLzilambda18354[147:140]};
  assign gzdLLzilambda15146 = {gzdLLzicase18351[7:0], gzdLLzicase18351[147:78], gzdLLzicase18351[77:8]};
  assign gzdLLzicase15143 = {gzdLLzilambda15146[139:70], gzdLLzilambda15146[147:140]};
  zdLLzicase15143  zdLLzicase15143 (gzdLLzicase15143[77:70], gzdLLzicase15143[69:62], gzdLLzicase15143[61:54], gzdLLzicase15143[53:46], gzdLLzicase15143[45:40], gzdLLzicase15143[39:23], gzdLLzicase15143[22:8], gzdLLzicase15143[7:0], callResR5);
  assign gzdLLzicase17968R1 = callResR5;
  zdLLzicase17968  zdLLzicase17968R1 (gzdLLzicase17968R1[69:0], callResR6);
  assign res = callResR6;
endmodule

module zdLLzicase17885 (input logic [69:0] arg0,
  input logic [16:0] arg1,
  output logic [143:0] res);
  logic [86:0] gzdLLzilambda14978;
  logic [139:0] gzdLLzilambda18120;
  logic [139:0] gzdLLzicase18021;
  logic [143:0] callRes;
  logic [160:0] gzdLLzilambda18115;
  logic [160:0] gzdLLzicase18112;
  logic [156:0] gzdLLzilambda14976;
  logic [86:0] gzdLLzicase14973;
  logic [69:0] callResR1;
  logic [69:0] gzdLLzicase17968;
  logic [143:0] callResR2;
  assign gzdLLzilambda14978 = {arg1, arg0};
  assign gzdLLzilambda18120 = {gzdLLzilambda14978[69:0], gzdLLzilambda14978[69:0]};
  assign gzdLLzicase18021 = gzdLLzilambda18120[139:0];
  zdLLzicase18021  zdLLzicase18021 (gzdLLzicase18021[139:70], gzdLLzicase18021[69:0], callRes);
  assign gzdLLzilambda18115 = {gzdLLzilambda14978[86:70], callRes};
  assign gzdLLzicase18112 = {gzdLLzilambda18115[143:0], gzdLLzilambda18115[160:144]};
  assign gzdLLzilambda14976 = {gzdLLzicase18112[16:0], gzdLLzicase18112[156:87], gzdLLzicase18112[86:17]};
  assign gzdLLzicase14973 = {gzdLLzilambda14976[139:70], gzdLLzilambda14976[156:140]};
  zdLLzicase14973  zdLLzicase14973 (gzdLLzicase14973[86:79], gzdLLzicase14973[78:71], gzdLLzicase14973[70:63], gzdLLzicase14973[62:55], gzdLLzicase14973[54:49], gzdLLzicase14973[48:32], gzdLLzicase14973[31:17], gzdLLzicase14973[16:0], callResR1);
  assign gzdLLzicase17968 = callResR1;
  zdLLzicase17968  zdLLzicase17968 (gzdLLzicase17968[69:0], callResR2);
  assign res = callResR2;
endmodule

module zdLLzicase17888 (input logic [7:0] arg0,
  input logic [69:0] arg1,
  output logic [143:0] res);
  assign res = {{4'h1, {6'h3e{1'h0}}}, arg0, arg1};
endmodule

module zdLLzicase17968 (input logic [69:0] arg0,
  output logic [143:0] res);
  assign res = {{3'h1, {7'h47{1'h0}}}, arg0};
endmodule

module zdLLzicase18021 (input logic [69:0] arg0,
  input logic [69:0] arg1,
  output logic [143:0] res);
  assign res = {4'h6, arg0, arg1};
endmodule

module zdLLzicase19243 (input logic [69:0] arg0,
  output logic [143:0] res);
  logic [69:0] gMainziloop;
  logic [139:0] gzdLLzilambda19507;
  logic [139:0] gzdLLzicase18021;
  logic [143:0] callRes;
  logic [143:0] gzdLLzilambda19502;
  logic [143:0] gzdLLzicase19500;
  logic [139:0] gzdLLzilambda15755;
  logic [69:0] gMainziinputs;
  logic [16:0] callResR1;
  logic [143:0] gzdLLzilambda19283;
  logic [143:0] gzdLLzicase19281;
  logic [86:0] gzdLLzilambda15753;
  logic [16:0] gMainziinstrIn;
  logic [16:0] gzdLLzicase14725;
  logic [143:0] gzdLLzilambda19278;
  logic [143:0] gzdLLzicase19276;
  logic [78:0] gzdLLzilambda15751;
  logic [139:0] gzdLLzilambda19273;
  logic [139:0] gzdLLzicase18021R1;
  logic [143:0] callResR2;
  logic [152:0] gzdLLzilambda19268;
  logic [152:0] gzdLLzicase19265;
  logic [148:0] gzdLLzilambda15749;
  logic [78:0] gzdLLzicase15735;
  logic [75:0] gzdLLzilambda15733;
  logic [139:0] gzdLLzilambda19240;
  logic [139:0] gzdLLzilambda15200;
  logic [77:0] callResR3;
  logic [77:0] gzdLLzilambda19235;
  logic [77:0] gzdLLzicase17888;
  logic [143:0] callResR4;
  logic [149:0] gzdLLzilambda19230;
  logic [149:0] gzdLLzicase19227;
  logic [83:0] gzdLLzilambda15731;
  logic [15:0] binOp;
  logic [15:0] binOpR1;
  logic [76:0] gzdLLzicase15648;
  logic [75:0] gzdLLzilambda15646;
  logic [139:0] gzdLLzilambda19088;
  logic [139:0] gzdLLzicase18021R2;
  logic [143:0] callResR5;
  logic [149:0] gzdLLzilambda19083;
  logic [149:0] gzdLLzicase19080;
  logic [145:0] gzdLLzilambda15644;
  logic [75:0] gzdLLzicase14914;
  logic [69:0] callResR6;
  logic [69:0] gzdLLzicase17968;
  logic [143:0] callResR7;
  logic [70:0] gzdLLzicase19223;
  logic [69:0] gzdLLzicase15649;
  logic [139:0] gzdLLzilambda18023;
  logic [139:0] gzdLLzicase18021R3;
  logic [143:0] callResR8;
  logic [143:0] gzdLLzilambda18018;
  logic [143:0] gzdLLzicase18016;
  logic [139:0] gzdLLzilambda15632;
  logic [69:0] gMainzipc;
  logic [5:0] callResR9;
  logic [143:0] gzdLLzilambda19071;
  logic [143:0] gzdLLzicase19069;
  logic [75:0] gzdLLzilambda15630;
  logic [11:0] binOpR2;
  logic [75:0] gzdLLzilambda15628;
  logic [139:0] gzdLLzilambda19066;
  logic [139:0] gzdLLzicase18021R4;
  logic [143:0] callResR10;
  logic [149:0] gzdLLzilambda19061;
  logic [149:0] gzdLLzicase19058;
  logic [145:0] gzdLLzilambda15626;
  logic [75:0] gzdLLzicase14914R1;
  logic [69:0] callResR11;
  logic [69:0] gzdLLzicase17968R1;
  logic [143:0] callResR12;
  logic [143:0] gzdLLzilambda19218;
  logic [143:0] gzdLLzicase19216;
  logic [69:0] gzdLLzilambda15728;
  logic [139:0] gzdLLzilambda19213;
  logic [139:0] gzdLLzicase18021R5;
  logic [143:0] callResR13;
  logic [143:0] gzdLLzilambda19208;
  logic [143:0] gzdLLzicase19206;
  logic [139:0] gzdLLzilambda15726;
  logic [69:0] gMainzipcR1;
  logic [5:0] callResR14;
  logic [143:0] gzdLLzilambda19203;
  logic [143:0] gzdLLzicase19201;
  logic [75:0] gzdLLzilambda15724;
  logic [75:0] gzdLLzilambda15676;
  logic [139:0] gzdLLzilambda19124;
  logic [139:0] gzdLLzicase18021R6;
  logic [143:0] callResR15;
  logic [149:0] gzdLLzilambda19119;
  logic [149:0] gzdLLzicase19116;
  logic [145:0] gzdLLzilambda15674;
  logic [69:0] gMainzioutputs;
  logic [14:0] callResR16;
  logic [149:0] gzdLLzilambda19112;
  logic [149:0] gzdLLzicase19109;
  logic [90:0] gzdLLzilambda15671;
  logic [20:0] gzdLLzicase14938;
  logic [14:0] callResR17;
  logic [84:0] gzdLLzilambda15663;
  logic [139:0] gzdLLzilambda19105;
  logic [139:0] gzdLLzicase18021R7;
  logic [143:0] callResR18;
  logic [158:0] gzdLLzilambda19100;
  logic [158:0] gzdLLzicase19097;
  logic [154:0] gzdLLzilambda15661;
  logic [84:0] gzdLLzicase14928;
  logic [69:0] callResR19;
  logic [69:0] gzdLLzicase17968R2;
  logic [143:0] callResR20;
  logic [143:0] gzdLLzilambda19198;
  logic [143:0] gzdLLzicase19196;
  logic [69:0] gzdLLzilambda15722;
  logic [139:0] gzdLLzilambda19193;
  logic [139:0] gzdLLzicase18021R8;
  logic [143:0] callResR21;
  logic [143:0] gzdLLzilambda19188;
  logic [143:0] gzdLLzicase19186;
  logic [139:0] gzdLLzilambda15720;
  logic [69:0] gMainzioutputsR1;
  logic [14:0] callResR22;
  logic [143:0] gzdLLzilambda19183;
  logic [143:0] gzdLLzicase19181;
  logic [84:0] gzdLLzilambda15718;
  logic [14:0] gzdLLzicase14964;
  logic [14:0] callResR23;
  logic [84:0] gzdLLzilambda15690;
  logic [139:0] gzdLLzilambda19141;
  logic [139:0] gzdLLzicase18021R9;
  logic [143:0] callResR24;
  logic [158:0] gzdLLzilambda19136;
  logic [158:0] gzdLLzicase19133;
  logic [154:0] gzdLLzilambda15688;
  logic [84:0] gzdLLzicase14928R1;
  logic [69:0] callResR25;
  logic [69:0] gzdLLzicase17968R3;
  logic [143:0] callResR26;
  logic [143:0] gzdLLzilambda19178;
  logic [143:0] gzdLLzicase19176;
  logic [69:0] gzdLLzilambda15716;
  logic [139:0] gzdLLzilambda19173;
  logic [139:0] gzdLLzicase18021R10;
  logic [143:0] callResR27;
  logic [143:0] gzdLLzilambda19168;
  logic [143:0] gzdLLzicase19166;
  logic [139:0] gzdLLzilambda15714;
  logic [69:0] gMainzioutputsR2;
  logic [14:0] callResR28;
  logic [143:0] gzdLLzilambda19163;
  logic [143:0] gzdLLzicase19161;
  logic [84:0] gzdLLzilambda15712;
  logic [78:0] gzdLLzicase15739;
  logic [75:0] gzdLLzilambda15612;
  logic [143:0] gzdLLzilambda15610;
  logic [143:0] gzdLLzilambda15607;
  logic [71:0] gzdLLzilambda15421;
  logic [71:0] gzdLLzicase18838;
  logic [69:0] gzdLLzicase15416;
  logic [139:0] gzdLLzilambda17895;
  logic [139:0] gzdLLzilambda15415;
  logic [77:0] callResR29;
  logic [77:0] gzdLLzilambda17890;
  logic [77:0] gzdLLzicase17888R1;
  logic [143:0] callResR30;
  logic [71:0] gzdLLzicase18840;
  logic [69:0] gzdLLzicase15417;
  logic [139:0] gzdLLzilambda17905;
  logic [139:0] gzdLLzilambda15413;
  logic [77:0] callResR31;
  logic [77:0] gzdLLzilambda17900;
  logic [77:0] gzdLLzicase17888R2;
  logic [143:0] callResR32;
  logic [71:0] gzdLLzicase18842;
  logic [69:0] gzdLLzicase15418;
  logic [139:0] gzdLLzilambda17915;
  logic [139:0] gzdLLzilambda15411;
  logic [77:0] callResR33;
  logic [77:0] gzdLLzilambda17910;
  logic [77:0] gzdLLzicase17888R3;
  logic [143:0] callResR34;
  logic [71:0] gzdLLzicase18844;
  logic [69:0] gzdLLzicase15419;
  logic [139:0] gzdLLzilambda17925;
  logic [139:0] gzdLLzilambda15200R1;
  logic [77:0] callResR35;
  logic [77:0] gzdLLzilambda17920;
  logic [77:0] gzdLLzicase17888R4;
  logic [143:0] callResR36;
  logic [147:0] gzdLLzilambda19049;
  logic [147:0] gzdLLzicase19045;
  logic [81:0] gzdLLzilambda15603;
  logic [71:0] gzdLLzilambda15435;
  logic [71:0] gzdLLzicase18846;
  logic [69:0] gzdLLzicase15430;
  logic [139:0] gzdLLzilambda17935;
  logic [139:0] gzdLLzilambda15415R1;
  logic [77:0] callResR37;
  logic [77:0] gzdLLzilambda17930;
  logic [77:0] gzdLLzicase17888R5;
  logic [143:0] callResR38;
  logic [71:0] gzdLLzicase18848;
  logic [69:0] gzdLLzicase15431;
  logic [139:0] gzdLLzilambda17945;
  logic [139:0] gzdLLzilambda15413R1;
  logic [77:0] callResR39;
  logic [77:0] gzdLLzilambda17940;
  logic [77:0] gzdLLzicase17888R6;
  logic [143:0] callResR40;
  logic [71:0] gzdLLzicase18850;
  logic [69:0] gzdLLzicase15432;
  logic [139:0] gzdLLzilambda17955;
  logic [139:0] gzdLLzilambda15411R1;
  logic [77:0] callResR41;
  logic [77:0] gzdLLzilambda17950;
  logic [77:0] gzdLLzicase17888R7;
  logic [143:0] callResR42;
  logic [71:0] gzdLLzicase18852;
  logic [69:0] gzdLLzicase15433;
  logic [139:0] gzdLLzilambda17965;
  logic [139:0] gzdLLzilambda15200R2;
  logic [77:0] callResR43;
  logic [77:0] gzdLLzilambda17960;
  logic [77:0] gzdLLzicase17888R8;
  logic [143:0] callResR44;
  logic [153:0] gzdLLzilambda19040;
  logic [153:0] gzdLLzicase19036;
  logic [87:0] gzdLLzilambda15599;
  logic [15:0] binOpR3;
  logic [7:0] unOp;
  logic [79:0] gzdLLzilambda15496;
  logic [141:0] gzdLLzilambda15494;
  logic [79:0] gzdLLzicase18855;
  logic [77:0] gzdLLzicase15485;
  logic [147:0] gzdLLzilambda17977;
  logic [147:0] gzdLLzicase17974;
  logic [147:0] gzdLLzilambda15483;
  logic [77:0] gzdLLzicase15480;
  logic [69:0] gzdLLzicase17968R4;
  logic [143:0] callResR45;
  logic [79:0] gzdLLzicase18858;
  logic [77:0] gzdLLzicase15487;
  logic [147:0] gzdLLzilambda17989;
  logic [147:0] gzdLLzicase17986;
  logic [147:0] gzdLLzilambda15471;
  logic [77:0] gzdLLzicase15468;
  logic [69:0] gzdLLzicase17968R5;
  logic [143:0] callResR46;
  logic [79:0] gzdLLzicase18861;
  logic [77:0] gzdLLzicase15489;
  logic [147:0] gzdLLzilambda18001;
  logic [147:0] gzdLLzicase17998;
  logic [147:0] gzdLLzilambda15459;
  logic [77:0] gzdLLzicase15456;
  logic [69:0] gzdLLzicase17968R6;
  logic [143:0] callResR47;
  logic [79:0] gzdLLzicase18864;
  logic [77:0] gzdLLzicase15491;
  logic [147:0] gzdLLzilambda18013;
  logic [147:0] gzdLLzicase18010;
  logic [147:0] gzdLLzilambda15447;
  logic [77:0] gzdLLzicase15143;
  logic [69:0] callResR48;
  logic [69:0] gzdLLzicase17968R7;
  logic [143:0] callResR49;
  logic [143:0] gzdLLzilambda19031;
  logic [143:0] gzdLLzicase19029;
  logic [69:0] gzdLLzilambda15595;
  logic [139:0] gzdLLzilambda19026;
  logic [139:0] gzdLLzicase18021R11;
  logic [143:0] callResR50;
  logic [143:0] gzdLLzilambda19021;
  logic [143:0] gzdLLzicase19019;
  logic [139:0] gzdLLzilambda15593;
  logic [69:0] gMainzipcR2;
  logic [5:0] callResR51;
  logic [143:0] gzdLLzilambda19016;
  logic [143:0] gzdLLzicase19014;
  logic [75:0] gzdLLzilambda15591;
  logic [11:0] binOpR4;
  logic [75:0] gzdLLzilambda15510;
  logic [139:0] gzdLLzilambda18881;
  logic [139:0] gzdLLzicase18021R12;
  logic [143:0] callResR52;
  logic [149:0] gzdLLzilambda18876;
  logic [149:0] gzdLLzicase18873;
  logic [145:0] gzdLLzilambda15508;
  logic [75:0] gzdLLzicase14914R2;
  logic [69:0] callResR53;
  logic [69:0] gzdLLzicase17968R8;
  logic [143:0] callResR54;
  logic [143:0] gzdLLzilambda19011;
  logic [143:0] gzdLLzicase19009;
  logic [69:0] gzdLLzilambda15589;
  logic [139:0] gzdLLzilambda19006;
  logic [139:0] gzdLLzicase18021R13;
  logic [143:0] callResR55;
  logic [143:0] gzdLLzilambda19001;
  logic [143:0] gzdLLzicase18999;
  logic [139:0] gzdLLzilambda15587;
  logic [69:0] gMainzipcR3;
  logic [5:0] callResR56;
  logic [143:0] gzdLLzilambda18996;
  logic [143:0] gzdLLzicase18994;
  logic [75:0] gzdLLzilambda15585;
  logic [75:0] gzdLLzilambda15537;
  logic [139:0] gzdLLzilambda18917;
  logic [139:0] gzdLLzicase18021R14;
  logic [143:0] callResR57;
  logic [149:0] gzdLLzilambda18912;
  logic [149:0] gzdLLzicase18909;
  logic [145:0] gzdLLzilambda15535;
  logic [69:0] gMainzioutputsR3;
  logic [14:0] callResR58;
  logic [149:0] gzdLLzilambda18905;
  logic [149:0] gzdLLzicase18902;
  logic [90:0] gzdLLzilambda15532;
  logic [20:0] gzdLLzicase14938R1;
  logic [14:0] callResR59;
  logic [84:0] gzdLLzilambda15524;
  logic [139:0] gzdLLzilambda18898;
  logic [139:0] gzdLLzicase18021R15;
  logic [143:0] callResR60;
  logic [158:0] gzdLLzilambda18893;
  logic [158:0] gzdLLzicase18890;
  logic [154:0] gzdLLzilambda15522;
  logic [84:0] gzdLLzicase14928R2;
  logic [69:0] callResR61;
  logic [69:0] gzdLLzicase17968R9;
  logic [143:0] callResR62;
  logic [143:0] gzdLLzilambda18991;
  logic [143:0] gzdLLzicase18989;
  logic [69:0] gzdLLzilambda15583;
  logic [139:0] gzdLLzilambda18986;
  logic [139:0] gzdLLzicase18021R16;
  logic [143:0] callResR63;
  logic [143:0] gzdLLzilambda18981;
  logic [143:0] gzdLLzicase18979;
  logic [139:0] gzdLLzilambda15581;
  logic [69:0] gMainzioutputsR4;
  logic [14:0] callResR64;
  logic [143:0] gzdLLzilambda18976;
  logic [143:0] gzdLLzicase18974;
  logic [84:0] gzdLLzilambda15579;
  logic [14:0] gzdLLzicase14964R1;
  logic [14:0] callResR65;
  logic [84:0] gzdLLzilambda15551;
  logic [139:0] gzdLLzilambda18934;
  logic [139:0] gzdLLzicase18021R17;
  logic [143:0] callResR66;
  logic [158:0] gzdLLzilambda18929;
  logic [158:0] gzdLLzicase18926;
  logic [154:0] gzdLLzilambda15549;
  logic [84:0] gzdLLzicase14928R3;
  logic [69:0] callResR67;
  logic [69:0] gzdLLzicase17968R10;
  logic [143:0] callResR68;
  logic [143:0] gzdLLzilambda18971;
  logic [143:0] gzdLLzicase18969;
  logic [69:0] gzdLLzilambda15577;
  logic [139:0] gzdLLzilambda18966;
  logic [139:0] gzdLLzicase18021R18;
  logic [143:0] callResR69;
  logic [143:0] gzdLLzilambda18961;
  logic [143:0] gzdLLzicase18959;
  logic [139:0] gzdLLzilambda15575;
  logic [69:0] gMainzioutputsR5;
  logic [14:0] callResR70;
  logic [143:0] gzdLLzilambda18956;
  logic [143:0] gzdLLzicase18954;
  logic [84:0] gzdLLzilambda15573;
  logic [78:0] gzdLLzicase15741;
  logic [75:0] gzdLLzilambda15407;
  logic [139:0] gzdLLzilambda18836;
  logic [139:0] gzdLLzilambda15200R3;
  logic [77:0] callResR71;
  logic [77:0] gzdLLzilambda18831;
  logic [77:0] gzdLLzicase17888R9;
  logic [143:0] callResR72;
  logic [149:0] gzdLLzilambda18826;
  logic [149:0] gzdLLzicase18823;
  logic [83:0] gzdLLzilambda15405;
  logic [75:0] gzdLLzilambda15227;
  logic [139:0] gzdLLzilambda18535;
  logic [139:0] gzdLLzicase18021R19;
  logic [143:0] callResR73;
  logic [149:0] gzdLLzilambda18530;
  logic [149:0] gzdLLzicase18527;
  logic [145:0] gzdLLzilambda15225;
  logic [69:0] gMainzioutputsR6;
  logic [14:0] callResR74;
  logic [149:0] gzdLLzilambda18523;
  logic [149:0] gzdLLzicase18520;
  logic [90:0] gzdLLzilambda15222;
  logic [20:0] gzdLLzicase14938R2;
  logic [14:0] callResR75;
  logic [84:0] gzdLLzilambda15214;
  logic [139:0] gzdLLzilambda18516;
  logic [139:0] gzdLLzicase18021R20;
  logic [143:0] callResR76;
  logic [158:0] gzdLLzilambda18511;
  logic [158:0] gzdLLzicase18508;
  logic [154:0] gzdLLzilambda15212;
  logic [84:0] gzdLLzicase14928R4;
  logic [69:0] callResR77;
  logic [69:0] gzdLLzicase17968R11;
  logic [143:0] callResR78;
  logic [151:0] gzdLLzilambda18819;
  logic [151:0] gzdLLzicase18816;
  logic [77:0] gzdLLzilambda15402;
  logic [77:0] gzdLLzilambda15254;
  logic [139:0] gzdLLzilambda18571;
  logic [139:0] gzdLLzicase18021R21;
  logic [143:0] callResR79;
  logic [151:0] gzdLLzilambda18566;
  logic [151:0] gzdLLzicase18563;
  logic [147:0] gzdLLzilambda15252;
  logic [69:0] gMainzioutputsR7;
  logic [14:0] callResR80;
  logic [151:0] gzdLLzilambda18559;
  logic [151:0] gzdLLzicase18556;
  logic [92:0] gzdLLzilambda15249;
  logic [22:0] gzdLLzicase15246;
  logic [84:0] gzdLLzilambda15241;
  logic [139:0] gzdLLzilambda18552;
  logic [139:0] gzdLLzicase18021R22;
  logic [143:0] callResR81;
  logic [158:0] gzdLLzilambda18547;
  logic [158:0] gzdLLzicase18544;
  logic [154:0] gzdLLzilambda15239;
  logic [84:0] gzdLLzicase14928R5;
  logic [69:0] callResR82;
  logic [69:0] gzdLLzicase17968R12;
  logic [143:0] callResR83;
  logic [143:0] gzdLLzilambda18812;
  logic [143:0] gzdLLzicase18810;
  logic [69:0] gzdLLzilambda15399;
  logic [139:0] gzdLLzilambda18807;
  logic [139:0] gzdLLzicase18021R23;
  logic [143:0] callResR84;
  logic [143:0] gzdLLzilambda18802;
  logic [143:0] gzdLLzicase18800;
  logic [139:0] gzdLLzilambda15397;
  logic [69:0] gMainzioutputsR8;
  logic [14:0] callResR85;
  logic [143:0] gzdLLzilambda18797;
  logic [143:0] gzdLLzicase18795;
  logic [84:0] gzdLLzilambda15395;
  logic [14:0] gzdLLzicase15272;
  logic [84:0] gzdLLzilambda15268;
  logic [139:0] gzdLLzilambda18588;
  logic [139:0] gzdLLzicase18021R24;
  logic [143:0] callResR86;
  logic [158:0] gzdLLzilambda18583;
  logic [158:0] gzdLLzicase18580;
  logic [154:0] gzdLLzilambda15266;
  logic [84:0] gzdLLzicase14928R6;
  logic [69:0] callResR87;
  logic [69:0] gzdLLzicase17968R13;
  logic [143:0] callResR88;
  logic [143:0] gzdLLzilambda18792;
  logic [143:0] gzdLLzicase18790;
  logic [69:0] gzdLLzilambda15393;
  logic [139:0] gzdLLzilambda18787;
  logic [139:0] gzdLLzicase18021R25;
  logic [143:0] callResR89;
  logic [143:0] gzdLLzilambda18782;
  logic [143:0] gzdLLzicase18780;
  logic [139:0] gzdLLzilambda15391;
  logic [69:0] gMainzioutputsR9;
  logic [14:0] callResR90;
  logic [143:0] gzdLLzilambda18777;
  logic [143:0] gzdLLzicase18775;
  logic [84:0] gzdLLzilambda15389;
  logic [78:0] gzdLLzicase15743;
  logic [75:0] gzdLLzilambda15198;
  logic [75:0] gzdLLzilambda15029;
  logic [139:0] gzdLLzilambda18221;
  logic [139:0] gzdLLzicase18021R26;
  logic [143:0] callResR91;
  logic [149:0] gzdLLzilambda18216;
  logic [149:0] gzdLLzicase18213;
  logic [145:0] gzdLLzilambda15027;
  logic [69:0] gMainzioutputsR10;
  logic [14:0] callResR92;
  logic [149:0] gzdLLzilambda18209;
  logic [149:0] gzdLLzicase18206;
  logic [90:0] gzdLLzilambda15024;
  logic [20:0] gzdLLzicase14938R3;
  logic [14:0] callResR93;
  logic [84:0] gzdLLzilambda15016;
  logic [139:0] gzdLLzilambda18202;
  logic [139:0] gzdLLzicase18021R27;
  logic [143:0] callResR94;
  logic [158:0] gzdLLzilambda18197;
  logic [158:0] gzdLLzicase18194;
  logic [154:0] gzdLLzilambda15014;
  logic [84:0] gzdLLzicase14928R7;
  logic [69:0] callResR95;
  logic [69:0] gzdLLzicase17968R14;
  logic [143:0] callResR96;
  logic [143:0] gzdLLzilambda18499;
  logic [143:0] gzdLLzicase18497;
  logic [69:0] gzdLLzilambda15196;
  logic [139:0] gzdLLzilambda18494;
  logic [139:0] gzdLLzicase18021R28;
  logic [143:0] callResR97;
  logic [143:0] gzdLLzilambda18489;
  logic [143:0] gzdLLzicase18487;
  logic [139:0] gzdLLzilambda15194;
  logic [69:0] gMainzioutputsR11;
  logic [14:0] callResR98;
  logic [143:0] gzdLLzilambda18484;
  logic [143:0] gzdLLzicase18482;
  logic [84:0] gzdLLzilambda15192;
  logic [14:0] gzdLLzicase14964R2;
  logic [14:0] callResR99;
  logic [84:0] gzdLLzilambda15043;
  logic [139:0] gzdLLzilambda18238;
  logic [139:0] gzdLLzicase18021R29;
  logic [143:0] callResR100;
  logic [158:0] gzdLLzilambda18233;
  logic [158:0] gzdLLzicase18230;
  logic [154:0] gzdLLzilambda15041;
  logic [84:0] gzdLLzicase14928R8;
  logic [69:0] callResR101;
  logic [69:0] gzdLLzicase17968R15;
  logic [143:0] callResR102;
  logic [143:0] gzdLLzilambda18479;
  logic [143:0] gzdLLzicase18477;
  logic [69:0] gzdLLzilambda15190;
  logic [139:0] gzdLLzilambda18474;
  logic [139:0] gzdLLzicase18021R30;
  logic [143:0] callResR103;
  logic [143:0] gzdLLzilambda18469;
  logic [143:0] gzdLLzicase18467;
  logic [139:0] gzdLLzilambda15188;
  logic [69:0] gMainzioutputsR12;
  logic [14:0] callResR104;
  logic [143:0] gzdLLzilambda18464;
  logic [143:0] gzdLLzicase18462;
  logic [84:0] gzdLLzilambda15186;
  logic [78:0] gzdLLzicase19261;
  logic [69:0] gzdLLzicase15744;
  logic [139:0] gzdLLzilambda18033;
  logic [139:0] gzdLLzicase18021R31;
  logic [143:0] callResR105;
  logic [143:0] gzdLLzilambda18028;
  logic [143:0] gzdLLzicase18026;
  logic [139:0] gzdLLzilambda15002;
  logic [69:0] gMainzipcR4;
  logic [5:0] callResR106;
  logic [143:0] gzdLLzilambda18185;
  logic [143:0] gzdLLzicase18183;
  logic [75:0] gzdLLzilambda15000;
  logic [11:0] binOpR5;
  logic [75:0] gzdLLzilambda14919;
  logic [139:0] gzdLLzilambda18050;
  logic [139:0] gzdLLzicase18021R32;
  logic [143:0] callResR107;
  logic [149:0] gzdLLzilambda18045;
  logic [149:0] gzdLLzicase18042;
  logic [145:0] gzdLLzilambda14917;
  logic [75:0] gzdLLzicase14914R3;
  logic [69:0] callResR108;
  logic [69:0] gzdLLzicase17968R16;
  logic [143:0] callResR109;
  logic [143:0] gzdLLzilambda18180;
  logic [143:0] gzdLLzicase18178;
  logic [69:0] gzdLLzilambda14998;
  logic [139:0] gzdLLzilambda18175;
  logic [139:0] gzdLLzicase18021R33;
  logic [143:0] callResR110;
  logic [143:0] gzdLLzilambda18170;
  logic [143:0] gzdLLzicase18168;
  logic [139:0] gzdLLzilambda14996;
  logic [69:0] gMainzipcR5;
  logic [5:0] callResR111;
  logic [143:0] gzdLLzilambda18165;
  logic [143:0] gzdLLzicase18163;
  logic [75:0] gzdLLzilambda14994;
  logic [75:0] gzdLLzilambda14946;
  logic [139:0] gzdLLzilambda18086;
  logic [139:0] gzdLLzicase18021R34;
  logic [143:0] callResR112;
  logic [149:0] gzdLLzilambda18081;
  logic [149:0] gzdLLzicase18078;
  logic [145:0] gzdLLzilambda14944;
  logic [69:0] gMainzioutputsR13;
  logic [14:0] callResR113;
  logic [149:0] gzdLLzilambda18074;
  logic [149:0] gzdLLzicase18071;
  logic [90:0] gzdLLzilambda14941;
  logic [20:0] gzdLLzicase14938R4;
  logic [14:0] callResR114;
  logic [84:0] gzdLLzilambda14933;
  logic [139:0] gzdLLzilambda18067;
  logic [139:0] gzdLLzicase18021R35;
  logic [143:0] callResR115;
  logic [158:0] gzdLLzilambda18062;
  logic [158:0] gzdLLzicase18059;
  logic [154:0] gzdLLzilambda14931;
  logic [84:0] gzdLLzicase14928R9;
  logic [69:0] callResR116;
  logic [69:0] gzdLLzicase17968R17;
  logic [143:0] callResR117;
  logic [143:0] gzdLLzilambda18160;
  logic [143:0] gzdLLzicase18158;
  logic [69:0] gzdLLzilambda14992;
  logic [139:0] gzdLLzilambda18155;
  logic [139:0] gzdLLzicase18021R36;
  logic [143:0] callResR118;
  logic [143:0] gzdLLzilambda18150;
  logic [143:0] gzdLLzicase18148;
  logic [139:0] gzdLLzilambda14990;
  logic [69:0] gMainzioutputsR14;
  logic [14:0] callResR119;
  logic [143:0] gzdLLzilambda18145;
  logic [143:0] gzdLLzicase18143;
  logic [84:0] gzdLLzilambda14988;
  logic [14:0] gzdLLzicase14964R3;
  logic [14:0] callResR120;
  logic [84:0] gzdLLzilambda14960;
  logic [139:0] gzdLLzilambda18103;
  logic [139:0] gzdLLzicase18021R37;
  logic [143:0] callResR121;
  logic [158:0] gzdLLzilambda18098;
  logic [158:0] gzdLLzicase18095;
  logic [154:0] gzdLLzilambda14958;
  logic [84:0] gzdLLzicase14928R10;
  logic [69:0] callResR122;
  logic [69:0] gzdLLzicase17968R18;
  logic [143:0] callResR123;
  logic [143:0] gzdLLzilambda18140;
  logic [143:0] gzdLLzicase18138;
  logic [69:0] gzdLLzilambda14986;
  logic [139:0] gzdLLzilambda18135;
  logic [139:0] gzdLLzicase18021R38;
  logic [143:0] callResR124;
  logic [143:0] gzdLLzilambda18130;
  logic [143:0] gzdLLzicase18128;
  logic [139:0] gzdLLzilambda14984;
  logic [69:0] gMainzioutputsR15;
  logic [14:0] callResR125;
  logic [143:0] gzdLLzilambda18125;
  logic [143:0] gzdLLzicase18123;
  logic [84:0] gzdLLzilambda14982;
  logic [143:0] gzdLLzilambda19245;
  logic [143:0] gzdLLzicase19243;
  logic [143:0] callResR126;
  assign gMainziloop = arg0;
  assign gzdLLzilambda19507 = {gMainziloop[69:0], gMainziloop[69:0]};
  assign gzdLLzicase18021 = gzdLLzilambda19507[139:0];
  zdLLzicase18021  zdLLzicase18021 (gzdLLzicase18021[139:70], gzdLLzicase18021[69:0], callRes);
  assign gzdLLzilambda19502 = callRes;
  assign gzdLLzicase19500 = gzdLLzilambda19502[143:0];
  assign gzdLLzilambda15755 = {gzdLLzicase19500[139:70], gzdLLzicase19500[69:0]};
  assign gMainziinputs = gzdLLzilambda15755[139:70];
  Mainziinputs  Mainziinputs (gMainziinputs[69:0], callResR1);
  assign gzdLLzilambda19283 = {{4'h3, {6'h35{1'h0}}}, callResR1, gzdLLzilambda15755[69:0]};
  assign gzdLLzicase19281 = gzdLLzilambda19283[143:0];
  assign gzdLLzilambda15753 = {gzdLLzicase19281[86:70], gzdLLzicase19281[69:0]};
  assign gMainziinstrIn = gzdLLzilambda15753[86:70];
  assign gzdLLzicase14725 = gMainziinstrIn[16:0];
  assign gzdLLzilambda19278 = {{2'h1, {6'h3f{1'h0}}}, gzdLLzicase14725[16:8], gzdLLzilambda15753[69:0]};
  assign gzdLLzicase19276 = gzdLLzilambda19278[143:0];
  assign gzdLLzilambda15751 = {gzdLLzicase19276[78:70], gzdLLzicase19276[69:0]};
  assign gzdLLzilambda19273 = {gzdLLzilambda15751[69:0], gzdLLzilambda15751[69:0]};
  assign gzdLLzicase18021R1 = gzdLLzilambda19273[139:0];
  zdLLzicase18021  zdLLzicase18021R1 (gzdLLzicase18021R1[139:70], gzdLLzicase18021R1[69:0], callResR2);
  assign gzdLLzilambda19268 = {gzdLLzilambda15751[78:70], callResR2};
  assign gzdLLzicase19265 = {gzdLLzilambda19268[143:0], gzdLLzilambda19268[152:144]};
  assign gzdLLzilambda15749 = {gzdLLzicase19265[8:0], gzdLLzicase19265[148:79], gzdLLzicase19265[78:9]};
  assign gzdLLzicase15735 = {gzdLLzilambda15749[148:140], gzdLLzilambda15749[69:0]};
  assign gzdLLzilambda15733 = {gzdLLzicase15735[75:70], gzdLLzicase15735[69:0]};
  assign gzdLLzilambda19240 = {gzdLLzilambda15733[69:0], gzdLLzilambda15733[69:0]};
  assign gzdLLzilambda15200 = gzdLLzilambda19240[139:0];
  zdLLzilambda15200  zdLLzilambda15200 (gzdLLzilambda15200[139:70], gzdLLzilambda15200[69:0], callResR3);
  assign gzdLLzilambda19235 = callResR3;
  assign gzdLLzicase17888 = gzdLLzilambda19235[77:0];
  zdLLzicase17888  zdLLzicase17888 (gzdLLzicase17888[77:70], gzdLLzicase17888[69:0], callResR4);
  assign gzdLLzilambda19230 = {gzdLLzilambda15733[75:70], callResR4};
  assign gzdLLzicase19227 = {gzdLLzilambda19230[143:0], gzdLLzilambda19230[149:144]};
  assign gzdLLzilambda15731 = {gzdLLzicase19227[5:0], gzdLLzicase19227[83:76], gzdLLzicase19227[75:6]};
  assign binOp = {gzdLLzilambda15731[77:70], 8'h00};
  assign binOpR1 = {gzdLLzilambda15731[77:70], 8'h00};
  assign gzdLLzicase15648 = {binOpR1[15:8] == binOpR1[7:0], gzdLLzilambda15731[83:78], gzdLLzilambda15731[69:0]};
  assign gzdLLzilambda15646 = {gzdLLzicase15648[75:70], gzdLLzicase15648[69:0]};
  assign gzdLLzilambda19088 = {gzdLLzilambda15646[69:0], gzdLLzilambda15646[69:0]};
  assign gzdLLzicase18021R2 = gzdLLzilambda19088[139:0];
  zdLLzicase18021  zdLLzicase18021R2 (gzdLLzicase18021R2[139:70], gzdLLzicase18021R2[69:0], callResR5);
  assign gzdLLzilambda19083 = {gzdLLzilambda15646[75:70], callResR5};
  assign gzdLLzicase19080 = {gzdLLzilambda19083[143:0], gzdLLzilambda19083[149:144]};
  assign gzdLLzilambda15644 = {gzdLLzicase19080[5:0], gzdLLzicase19080[145:76], gzdLLzicase19080[75:6]};
  assign gzdLLzicase14914 = {gzdLLzilambda15644[139:70], gzdLLzilambda15644[145:140]};
  zdLLzicase14914  zdLLzicase14914 (gzdLLzicase14914[75:68], gzdLLzicase14914[67:60], gzdLLzicase14914[59:52], gzdLLzicase14914[51:44], gzdLLzicase14914[43:38], gzdLLzicase14914[37:21], gzdLLzicase14914[20:6], gzdLLzicase14914[5:0], callResR6);
  assign gzdLLzicase17968 = callResR6;
  zdLLzicase17968  zdLLzicase17968 (gzdLLzicase17968[69:0], callResR7);
  assign gzdLLzicase19223 = {binOp[15:8] == binOp[7:0], gzdLLzilambda15731[69:0]};
  assign gzdLLzicase15649 = gzdLLzicase19223[69:0];
  assign gzdLLzilambda18023 = {gzdLLzicase15649[69:0], gzdLLzicase15649[69:0]};
  assign gzdLLzicase18021R3 = gzdLLzilambda18023[139:0];
  zdLLzicase18021  zdLLzicase18021R3 (gzdLLzicase18021R3[139:70], gzdLLzicase18021R3[69:0], callResR8);
  assign gzdLLzilambda18018 = callResR8;
  assign gzdLLzicase18016 = gzdLLzilambda18018[143:0];
  assign gzdLLzilambda15632 = {gzdLLzicase18016[139:70], gzdLLzicase18016[69:0]};
  assign gMainzipc = gzdLLzilambda15632[139:70];
  Mainzipc  Mainzipc (gMainzipc[69:0], callResR9);
  assign gzdLLzilambda19071 = {{7'h44{1'h0}}, callResR9, gzdLLzilambda15632[69:0]};
  assign gzdLLzicase19069 = gzdLLzilambda19071[143:0];
  assign gzdLLzilambda15630 = {gzdLLzicase19069[75:70], gzdLLzicase19069[69:0]};
  assign binOpR2 = {gzdLLzilambda15630[75:70], 6'h01};
  assign gzdLLzilambda15628 = {binOpR2[11:6] + binOpR2[5:0], gzdLLzilambda15630[69:0]};
  assign gzdLLzilambda19066 = {gzdLLzilambda15628[69:0], gzdLLzilambda15628[69:0]};
  assign gzdLLzicase18021R4 = gzdLLzilambda19066[139:0];
  zdLLzicase18021  zdLLzicase18021R4 (gzdLLzicase18021R4[139:70], gzdLLzicase18021R4[69:0], callResR10);
  assign gzdLLzilambda19061 = {gzdLLzilambda15628[75:70], callResR10};
  assign gzdLLzicase19058 = {gzdLLzilambda19061[143:0], gzdLLzilambda19061[149:144]};
  assign gzdLLzilambda15626 = {gzdLLzicase19058[5:0], gzdLLzicase19058[145:76], gzdLLzicase19058[75:6]};
  assign gzdLLzicase14914R1 = {gzdLLzilambda15626[139:70], gzdLLzilambda15626[145:140]};
  zdLLzicase14914  zdLLzicase14914R1 (gzdLLzicase14914R1[75:68], gzdLLzicase14914R1[67:60], gzdLLzicase14914R1[59:52], gzdLLzicase14914R1[51:44], gzdLLzicase14914R1[43:38], gzdLLzicase14914R1[37:21], gzdLLzicase14914R1[20:6], gzdLLzicase14914R1[5:0], callResR11);
  assign gzdLLzicase17968R1 = callResR11;
  zdLLzicase17968  zdLLzicase17968R1 (gzdLLzicase17968R1[69:0], callResR12);
  assign gzdLLzilambda19218 = (gzdLLzicase19223[70] == 1'h1) ? callResR12 : callResR7;
  assign gzdLLzicase19216 = gzdLLzilambda19218[143:0];
  assign gzdLLzilambda15728 = gzdLLzicase19216[69:0];
  assign gzdLLzilambda19213 = {gzdLLzilambda15728[69:0], gzdLLzilambda15728[69:0]};
  assign gzdLLzicase18021R5 = gzdLLzilambda19213[139:0];
  zdLLzicase18021  zdLLzicase18021R5 (gzdLLzicase18021R5[139:70], gzdLLzicase18021R5[69:0], callResR13);
  assign gzdLLzilambda19208 = callResR13;
  assign gzdLLzicase19206 = gzdLLzilambda19208[143:0];
  assign gzdLLzilambda15726 = {gzdLLzicase19206[139:70], gzdLLzicase19206[69:0]};
  assign gMainzipcR1 = gzdLLzilambda15726[139:70];
  Mainzipc  MainzipcR1 (gMainzipcR1[69:0], callResR14);
  assign gzdLLzilambda19203 = {{7'h44{1'h0}}, callResR14, gzdLLzilambda15726[69:0]};
  assign gzdLLzicase19201 = gzdLLzilambda19203[143:0];
  assign gzdLLzilambda15724 = {gzdLLzicase19201[75:70], gzdLLzicase19201[69:0]};
  assign gzdLLzilambda15676 = {gzdLLzilambda15724[75:70], gzdLLzilambda15724[69:0]};
  assign gzdLLzilambda19124 = {gzdLLzilambda15676[69:0], gzdLLzilambda15676[69:0]};
  assign gzdLLzicase18021R6 = gzdLLzilambda19124[139:0];
  zdLLzicase18021  zdLLzicase18021R6 (gzdLLzicase18021R6[139:70], gzdLLzicase18021R6[69:0], callResR15);
  assign gzdLLzilambda19119 = {gzdLLzilambda15676[75:70], callResR15};
  assign gzdLLzicase19116 = {gzdLLzilambda19119[143:0], gzdLLzilambda19119[149:144]};
  assign gzdLLzilambda15674 = {gzdLLzicase19116[5:0], gzdLLzicase19116[145:76], gzdLLzicase19116[75:6]};
  assign gMainzioutputs = gzdLLzilambda15674[139:70];
  Mainzioutputs  Mainzioutputs (gMainzioutputs[69:0], callResR16);
  assign gzdLLzilambda19112 = {gzdLLzilambda15674[145:140], {4'h5, {6'h37{1'h0}}}, callResR16, gzdLLzilambda15674[69:0]};
  assign gzdLLzicase19109 = {gzdLLzilambda19112[143:0], gzdLLzilambda19112[149:144]};
  assign gzdLLzilambda15671 = {gzdLLzicase19109[5:0], gzdLLzicase19109[90:76], gzdLLzicase19109[75:6]};
  assign gzdLLzicase14938 = {gzdLLzilambda15671[84:70], gzdLLzilambda15671[90:85]};
  zdLLzicase14938  zdLLzicase14938 (gzdLLzicase14938[20], gzdLLzicase14938[19:14], gzdLLzicase14938[13:6], gzdLLzicase14938[5:0], callResR17);
  assign gzdLLzilambda15663 = {callResR17, gzdLLzilambda15671[69:0]};
  assign gzdLLzilambda19105 = {gzdLLzilambda15663[69:0], gzdLLzilambda15663[69:0]};
  assign gzdLLzicase18021R7 = gzdLLzilambda19105[139:0];
  zdLLzicase18021  zdLLzicase18021R7 (gzdLLzicase18021R7[139:70], gzdLLzicase18021R7[69:0], callResR18);
  assign gzdLLzilambda19100 = {gzdLLzilambda15663[84:70], callResR18};
  assign gzdLLzicase19097 = {gzdLLzilambda19100[143:0], gzdLLzilambda19100[158:144]};
  assign gzdLLzilambda15661 = {gzdLLzicase19097[14:0], gzdLLzicase19097[154:85], gzdLLzicase19097[84:15]};
  assign gzdLLzicase14928 = {gzdLLzilambda15661[139:70], gzdLLzilambda15661[154:140]};
  zdLLzicase14928  zdLLzicase14928 (gzdLLzicase14928[84:77], gzdLLzicase14928[76:69], gzdLLzicase14928[68:61], gzdLLzicase14928[60:53], gzdLLzicase14928[52:47], gzdLLzicase14928[46:30], gzdLLzicase14928[29:15], gzdLLzicase14928[14:0], callResR19);
  assign gzdLLzicase17968R2 = callResR19;
  zdLLzicase17968  zdLLzicase17968R2 (gzdLLzicase17968R2[69:0], callResR20);
  assign gzdLLzilambda19198 = callResR20;
  assign gzdLLzicase19196 = gzdLLzilambda19198[143:0];
  assign gzdLLzilambda15722 = gzdLLzicase19196[69:0];
  assign gzdLLzilambda19193 = {gzdLLzilambda15722[69:0], gzdLLzilambda15722[69:0]};
  assign gzdLLzicase18021R8 = gzdLLzilambda19193[139:0];
  zdLLzicase18021  zdLLzicase18021R8 (gzdLLzicase18021R8[139:70], gzdLLzicase18021R8[69:0], callResR21);
  assign gzdLLzilambda19188 = callResR21;
  assign gzdLLzicase19186 = gzdLLzilambda19188[143:0];
  assign gzdLLzilambda15720 = {gzdLLzicase19186[139:70], gzdLLzicase19186[69:0]};
  assign gMainzioutputsR1 = gzdLLzilambda15720[139:70];
  Mainzioutputs  MainzioutputsR1 (gMainzioutputsR1[69:0], callResR22);
  assign gzdLLzilambda19183 = {{4'h5, {6'h37{1'h0}}}, callResR22, gzdLLzilambda15720[69:0]};
  assign gzdLLzicase19181 = gzdLLzilambda19183[143:0];
  assign gzdLLzilambda15718 = {gzdLLzicase19181[84:70], gzdLLzicase19181[69:0]};
  assign gzdLLzicase14964 = gzdLLzilambda15718[84:70];
  zdLLzicase14964  zdLLzicase14964 (gzdLLzicase14964[14], gzdLLzicase14964[13:8], gzdLLzicase14964[7:0], callResR23);
  assign gzdLLzilambda15690 = {callResR23, gzdLLzilambda15718[69:0]};
  assign gzdLLzilambda19141 = {gzdLLzilambda15690[69:0], gzdLLzilambda15690[69:0]};
  assign gzdLLzicase18021R9 = gzdLLzilambda19141[139:0];
  zdLLzicase18021  zdLLzicase18021R9 (gzdLLzicase18021R9[139:70], gzdLLzicase18021R9[69:0], callResR24);
  assign gzdLLzilambda19136 = {gzdLLzilambda15690[84:70], callResR24};
  assign gzdLLzicase19133 = {gzdLLzilambda19136[143:0], gzdLLzilambda19136[158:144]};
  assign gzdLLzilambda15688 = {gzdLLzicase19133[14:0], gzdLLzicase19133[154:85], gzdLLzicase19133[84:15]};
  assign gzdLLzicase14928R1 = {gzdLLzilambda15688[139:70], gzdLLzilambda15688[154:140]};
  zdLLzicase14928  zdLLzicase14928R1 (gzdLLzicase14928R1[84:77], gzdLLzicase14928R1[76:69], gzdLLzicase14928R1[68:61], gzdLLzicase14928R1[60:53], gzdLLzicase14928R1[52:47], gzdLLzicase14928R1[46:30], gzdLLzicase14928R1[29:15], gzdLLzicase14928R1[14:0], callResR25);
  assign gzdLLzicase17968R3 = callResR25;
  zdLLzicase17968  zdLLzicase17968R3 (gzdLLzicase17968R3[69:0], callResR26);
  assign gzdLLzilambda19178 = callResR26;
  assign gzdLLzicase19176 = gzdLLzilambda19178[143:0];
  assign gzdLLzilambda15716 = gzdLLzicase19176[69:0];
  assign gzdLLzilambda19173 = {gzdLLzilambda15716[69:0], gzdLLzilambda15716[69:0]};
  assign gzdLLzicase18021R10 = gzdLLzilambda19173[139:0];
  zdLLzicase18021  zdLLzicase18021R10 (gzdLLzicase18021R10[139:70], gzdLLzicase18021R10[69:0], callResR27);
  assign gzdLLzilambda19168 = callResR27;
  assign gzdLLzicase19166 = gzdLLzilambda19168[143:0];
  assign gzdLLzilambda15714 = {gzdLLzicase19166[139:70], gzdLLzicase19166[69:0]};
  assign gMainzioutputsR2 = gzdLLzilambda15714[139:70];
  Mainzioutputs  MainzioutputsR2 (gMainzioutputsR2[69:0], callResR28);
  assign gzdLLzilambda19163 = {{4'h5, {6'h37{1'h0}}}, callResR28, gzdLLzilambda15714[69:0]};
  assign gzdLLzicase19161 = gzdLLzilambda19163[143:0];
  assign gzdLLzilambda15712 = {gzdLLzicase19161[84:70], gzdLLzicase19161[69:0]};
  assign gzdLLzicase15739 = {gzdLLzilambda15749[148:140], gzdLLzilambda15749[69:0]};
  assign gzdLLzilambda15612 = {gzdLLzicase15739[75:74], gzdLLzicase15739[73:72], gzdLLzicase15739[71:70], gzdLLzicase15739[69:0]};
  assign gzdLLzilambda15610 = {gzdLLzilambda15612[75:74], gzdLLzilambda15612[73:72], gzdLLzilambda15612[71:70], gzdLLzilambda15612[69:0]};
  assign gzdLLzilambda15607 = {gzdLLzilambda15610[141:72], gzdLLzilambda15610[143:142], gzdLLzilambda15610[71:70], gzdLLzilambda15610[69:0]};
  assign gzdLLzilambda15421 = {gzdLLzilambda15607[143:142], gzdLLzilambda15607[69:0]};
  assign gzdLLzicase18838 = {gzdLLzilambda15421[71:70], gzdLLzilambda15421[69:0]};
  assign gzdLLzicase15416 = gzdLLzicase18838[69:0];
  assign gzdLLzilambda17895 = {gzdLLzicase15416[69:0], gzdLLzicase15416[69:0]};
  assign gzdLLzilambda15415 = gzdLLzilambda17895[139:0];
  zdLLzilambda15415  zdLLzilambda15415 (gzdLLzilambda15415[139:70], gzdLLzilambda15415[69:0], callResR29);
  assign gzdLLzilambda17890 = callResR29;
  assign gzdLLzicase17888R1 = gzdLLzilambda17890[77:0];
  zdLLzicase17888  zdLLzicase17888R1 (gzdLLzicase17888R1[77:70], gzdLLzicase17888R1[69:0], callResR30);
  assign gzdLLzicase18840 = {gzdLLzilambda15421[71:70], gzdLLzilambda15421[69:0]};
  assign gzdLLzicase15417 = gzdLLzicase18840[69:0];
  assign gzdLLzilambda17905 = {gzdLLzicase15417[69:0], gzdLLzicase15417[69:0]};
  assign gzdLLzilambda15413 = gzdLLzilambda17905[139:0];
  zdLLzilambda15413  zdLLzilambda15413 (gzdLLzilambda15413[139:70], gzdLLzilambda15413[69:0], callResR31);
  assign gzdLLzilambda17900 = callResR31;
  assign gzdLLzicase17888R2 = gzdLLzilambda17900[77:0];
  zdLLzicase17888  zdLLzicase17888R2 (gzdLLzicase17888R2[77:70], gzdLLzicase17888R2[69:0], callResR32);
  assign gzdLLzicase18842 = {gzdLLzilambda15421[71:70], gzdLLzilambda15421[69:0]};
  assign gzdLLzicase15418 = gzdLLzicase18842[69:0];
  assign gzdLLzilambda17915 = {gzdLLzicase15418[69:0], gzdLLzicase15418[69:0]};
  assign gzdLLzilambda15411 = gzdLLzilambda17915[139:0];
  zdLLzilambda15411  zdLLzilambda15411 (gzdLLzilambda15411[139:70], gzdLLzilambda15411[69:0], callResR33);
  assign gzdLLzilambda17910 = callResR33;
  assign gzdLLzicase17888R3 = gzdLLzilambda17910[77:0];
  zdLLzicase17888  zdLLzicase17888R3 (gzdLLzicase17888R3[77:70], gzdLLzicase17888R3[69:0], callResR34);
  assign gzdLLzicase18844 = {gzdLLzilambda15421[71:70], gzdLLzilambda15421[69:0]};
  assign gzdLLzicase15419 = gzdLLzicase18844[69:0];
  assign gzdLLzilambda17925 = {gzdLLzicase15419[69:0], gzdLLzicase15419[69:0]};
  assign gzdLLzilambda15200R1 = gzdLLzilambda17925[139:0];
  zdLLzilambda15200  zdLLzilambda15200R1 (gzdLLzilambda15200R1[139:70], gzdLLzilambda15200R1[69:0], callResR35);
  assign gzdLLzilambda17920 = callResR35;
  assign gzdLLzicase17888R4 = gzdLLzilambda17920[77:0];
  zdLLzicase17888  zdLLzicase17888R4 (gzdLLzicase17888R4[77:70], gzdLLzicase17888R4[69:0], callResR36);
  assign gzdLLzilambda19049 = {gzdLLzilambda15607[139:70], gzdLLzilambda15607[141:140], (gzdLLzicase18844[71:70] == 2'h0) ? callResR36 : ((gzdLLzicase18842[71:70] == 2'h1) ? callResR34 : ((gzdLLzicase18840[71:70] == 2'h2) ? callResR32 : callResR30))};
  assign gzdLLzicase19045 = {gzdLLzilambda19049[143:0], gzdLLzilambda19049[147:146], gzdLLzilambda19049[145:144]};
  assign gzdLLzilambda15603 = {gzdLLzicase19045[3:2], gzdLLzicase19045[1:0], gzdLLzicase19045[81:74], gzdLLzicase19045[73:4]};
  assign gzdLLzilambda15435 = {gzdLLzilambda15603[81:80], gzdLLzilambda15603[69:0]};
  assign gzdLLzicase18846 = {gzdLLzilambda15435[71:70], gzdLLzilambda15435[69:0]};
  assign gzdLLzicase15430 = gzdLLzicase18846[69:0];
  assign gzdLLzilambda17935 = {gzdLLzicase15430[69:0], gzdLLzicase15430[69:0]};
  assign gzdLLzilambda15415R1 = gzdLLzilambda17935[139:0];
  zdLLzilambda15415  zdLLzilambda15415R1 (gzdLLzilambda15415R1[139:70], gzdLLzilambda15415R1[69:0], callResR37);
  assign gzdLLzilambda17930 = callResR37;
  assign gzdLLzicase17888R5 = gzdLLzilambda17930[77:0];
  zdLLzicase17888  zdLLzicase17888R5 (gzdLLzicase17888R5[77:70], gzdLLzicase17888R5[69:0], callResR38);
  assign gzdLLzicase18848 = {gzdLLzilambda15435[71:70], gzdLLzilambda15435[69:0]};
  assign gzdLLzicase15431 = gzdLLzicase18848[69:0];
  assign gzdLLzilambda17945 = {gzdLLzicase15431[69:0], gzdLLzicase15431[69:0]};
  assign gzdLLzilambda15413R1 = gzdLLzilambda17945[139:0];
  zdLLzilambda15413  zdLLzilambda15413R1 (gzdLLzilambda15413R1[139:70], gzdLLzilambda15413R1[69:0], callResR39);
  assign gzdLLzilambda17940 = callResR39;
  assign gzdLLzicase17888R6 = gzdLLzilambda17940[77:0];
  zdLLzicase17888  zdLLzicase17888R6 (gzdLLzicase17888R6[77:70], gzdLLzicase17888R6[69:0], callResR40);
  assign gzdLLzicase18850 = {gzdLLzilambda15435[71:70], gzdLLzilambda15435[69:0]};
  assign gzdLLzicase15432 = gzdLLzicase18850[69:0];
  assign gzdLLzilambda17955 = {gzdLLzicase15432[69:0], gzdLLzicase15432[69:0]};
  assign gzdLLzilambda15411R1 = gzdLLzilambda17955[139:0];
  zdLLzilambda15411  zdLLzilambda15411R1 (gzdLLzilambda15411R1[139:70], gzdLLzilambda15411R1[69:0], callResR41);
  assign gzdLLzilambda17950 = callResR41;
  assign gzdLLzicase17888R7 = gzdLLzilambda17950[77:0];
  zdLLzicase17888  zdLLzicase17888R7 (gzdLLzicase17888R7[77:70], gzdLLzicase17888R7[69:0], callResR42);
  assign gzdLLzicase18852 = {gzdLLzilambda15435[71:70], gzdLLzilambda15435[69:0]};
  assign gzdLLzicase15433 = gzdLLzicase18852[69:0];
  assign gzdLLzilambda17965 = {gzdLLzicase15433[69:0], gzdLLzicase15433[69:0]};
  assign gzdLLzilambda15200R2 = gzdLLzilambda17965[139:0];
  zdLLzilambda15200  zdLLzilambda15200R2 (gzdLLzilambda15200R2[139:70], gzdLLzilambda15200R2[69:0], callResR43);
  assign gzdLLzilambda17960 = callResR43;
  assign gzdLLzicase17888R8 = gzdLLzilambda17960[77:0];
  zdLLzicase17888  zdLLzicase17888R8 (gzdLLzicase17888R8[77:70], gzdLLzicase17888R8[69:0], callResR44);
  assign gzdLLzilambda19040 = {gzdLLzilambda15603[79:78], gzdLLzilambda15603[77:70], (gzdLLzicase18852[71:70] == 2'h0) ? callResR44 : ((gzdLLzicase18850[71:70] == 2'h1) ? callResR42 : ((gzdLLzicase18848[71:70] == 2'h2) ? callResR40 : callResR38))};
  assign gzdLLzicase19036 = {gzdLLzilambda19040[143:0], gzdLLzilambda19040[153:152], gzdLLzilambda19040[151:144]};
  assign gzdLLzilambda15599 = {gzdLLzicase19036[9:8], gzdLLzicase19036[7:0], gzdLLzicase19036[87:80], gzdLLzicase19036[79:10]};
  assign binOpR3 = {gzdLLzilambda15599[85:78], gzdLLzilambda15599[77:70]};
  assign unOp = binOpR3[15:8] & binOpR3[7:0];
  assign gzdLLzilambda15496 = {gzdLLzilambda15599[87:86], ~unOp[7:0], gzdLLzilambda15599[69:0]};
  assign gzdLLzilambda15494 = {gzdLLzilambda15496[79:78], gzdLLzilambda15496[77:70], gzdLLzilambda15496[69:0]};
  assign gzdLLzicase18855 = {gzdLLzilambda15494[141:140], gzdLLzilambda15494[139:70], gzdLLzilambda15494[69:0]};
  assign gzdLLzicase15485 = {gzdLLzicase18855[77:70], gzdLLzicase18855[69:0]};
  assign gzdLLzilambda17977 = {gzdLLzicase15485[77:70], gzdLLzicase15485[69:0], gzdLLzicase15485[69:0]};
  assign gzdLLzicase17974 = {gzdLLzilambda17977[139:0], gzdLLzilambda17977[147:140]};
  assign gzdLLzilambda15483 = {gzdLLzicase17974[7:0], gzdLLzicase17974[147:78], gzdLLzicase17974[77:8]};
  assign gzdLLzicase15480 = {gzdLLzilambda15483[139:70], gzdLLzilambda15483[147:140]};
  assign gzdLLzicase17968R4 = {gzdLLzicase15480[77:70], gzdLLzicase15480[69:62], gzdLLzicase15480[61:54], gzdLLzicase15480[7:0], gzdLLzicase15480[45:40], gzdLLzicase15480[39:23], gzdLLzicase15480[22:8]};
  zdLLzicase17968  zdLLzicase17968R4 (gzdLLzicase17968R4[69:0], callResR45);
  assign gzdLLzicase18858 = {gzdLLzilambda15494[141:140], gzdLLzilambda15494[139:70], gzdLLzilambda15494[69:0]};
  assign gzdLLzicase15487 = {gzdLLzicase18858[77:70], gzdLLzicase18858[69:0]};
  assign gzdLLzilambda17989 = {gzdLLzicase15487[77:70], gzdLLzicase15487[69:0], gzdLLzicase15487[69:0]};
  assign gzdLLzicase17986 = {gzdLLzilambda17989[139:0], gzdLLzilambda17989[147:140]};
  assign gzdLLzilambda15471 = {gzdLLzicase17986[7:0], gzdLLzicase17986[147:78], gzdLLzicase17986[77:8]};
  assign gzdLLzicase15468 = {gzdLLzilambda15471[139:70], gzdLLzilambda15471[147:140]};
  assign gzdLLzicase17968R5 = {gzdLLzicase15468[77:70], gzdLLzicase15468[69:62], gzdLLzicase15468[7:0], gzdLLzicase15468[53:46], gzdLLzicase15468[45:40], gzdLLzicase15468[39:23], gzdLLzicase15468[22:8]};
  zdLLzicase17968  zdLLzicase17968R5 (gzdLLzicase17968R5[69:0], callResR46);
  assign gzdLLzicase18861 = {gzdLLzilambda15494[141:140], gzdLLzilambda15494[139:70], gzdLLzilambda15494[69:0]};
  assign gzdLLzicase15489 = {gzdLLzicase18861[77:70], gzdLLzicase18861[69:0]};
  assign gzdLLzilambda18001 = {gzdLLzicase15489[77:70], gzdLLzicase15489[69:0], gzdLLzicase15489[69:0]};
  assign gzdLLzicase17998 = {gzdLLzilambda18001[139:0], gzdLLzilambda18001[147:140]};
  assign gzdLLzilambda15459 = {gzdLLzicase17998[7:0], gzdLLzicase17998[147:78], gzdLLzicase17998[77:8]};
  assign gzdLLzicase15456 = {gzdLLzilambda15459[139:70], gzdLLzilambda15459[147:140]};
  assign gzdLLzicase17968R6 = {gzdLLzicase15456[77:70], gzdLLzicase15456[7:0], gzdLLzicase15456[61:54], gzdLLzicase15456[53:46], gzdLLzicase15456[45:40], gzdLLzicase15456[39:23], gzdLLzicase15456[22:8]};
  zdLLzicase17968  zdLLzicase17968R6 (gzdLLzicase17968R6[69:0], callResR47);
  assign gzdLLzicase18864 = {gzdLLzilambda15494[141:140], gzdLLzilambda15494[139:70], gzdLLzilambda15494[69:0]};
  assign gzdLLzicase15491 = {gzdLLzicase18864[77:70], gzdLLzicase18864[69:0]};
  assign gzdLLzilambda18013 = {gzdLLzicase15491[77:70], gzdLLzicase15491[69:0], gzdLLzicase15491[69:0]};
  assign gzdLLzicase18010 = {gzdLLzilambda18013[139:0], gzdLLzilambda18013[147:140]};
  assign gzdLLzilambda15447 = {gzdLLzicase18010[7:0], gzdLLzicase18010[147:78], gzdLLzicase18010[77:8]};
  assign gzdLLzicase15143 = {gzdLLzilambda15447[139:70], gzdLLzilambda15447[147:140]};
  zdLLzicase15143  zdLLzicase15143 (gzdLLzicase15143[77:70], gzdLLzicase15143[69:62], gzdLLzicase15143[61:54], gzdLLzicase15143[53:46], gzdLLzicase15143[45:40], gzdLLzicase15143[39:23], gzdLLzicase15143[22:8], gzdLLzicase15143[7:0], callResR48);
  assign gzdLLzicase17968R7 = callResR48;
  zdLLzicase17968  zdLLzicase17968R7 (gzdLLzicase17968R7[69:0], callResR49);
  assign gzdLLzilambda19031 = (gzdLLzicase18864[79:78] == 2'h0) ? callResR49 : ((gzdLLzicase18861[79:78] == 2'h1) ? callResR47 : ((gzdLLzicase18858[79:78] == 2'h2) ? callResR46 : callResR45));
  assign gzdLLzicase19029 = gzdLLzilambda19031[143:0];
  assign gzdLLzilambda15595 = gzdLLzicase19029[69:0];
  assign gzdLLzilambda19026 = {gzdLLzilambda15595[69:0], gzdLLzilambda15595[69:0]};
  assign gzdLLzicase18021R11 = gzdLLzilambda19026[139:0];
  zdLLzicase18021  zdLLzicase18021R11 (gzdLLzicase18021R11[139:70], gzdLLzicase18021R11[69:0], callResR50);
  assign gzdLLzilambda19021 = callResR50;
  assign gzdLLzicase19019 = gzdLLzilambda19021[143:0];
  assign gzdLLzilambda15593 = {gzdLLzicase19019[139:70], gzdLLzicase19019[69:0]};
  assign gMainzipcR2 = gzdLLzilambda15593[139:70];
  Mainzipc  MainzipcR2 (gMainzipcR2[69:0], callResR51);
  assign gzdLLzilambda19016 = {{7'h44{1'h0}}, callResR51, gzdLLzilambda15593[69:0]};
  assign gzdLLzicase19014 = gzdLLzilambda19016[143:0];
  assign gzdLLzilambda15591 = {gzdLLzicase19014[75:70], gzdLLzicase19014[69:0]};
  assign binOpR4 = {gzdLLzilambda15591[75:70], 6'h01};
  assign gzdLLzilambda15510 = {binOpR4[11:6] + binOpR4[5:0], gzdLLzilambda15591[69:0]};
  assign gzdLLzilambda18881 = {gzdLLzilambda15510[69:0], gzdLLzilambda15510[69:0]};
  assign gzdLLzicase18021R12 = gzdLLzilambda18881[139:0];
  zdLLzicase18021  zdLLzicase18021R12 (gzdLLzicase18021R12[139:70], gzdLLzicase18021R12[69:0], callResR52);
  assign gzdLLzilambda18876 = {gzdLLzilambda15510[75:70], callResR52};
  assign gzdLLzicase18873 = {gzdLLzilambda18876[143:0], gzdLLzilambda18876[149:144]};
  assign gzdLLzilambda15508 = {gzdLLzicase18873[5:0], gzdLLzicase18873[145:76], gzdLLzicase18873[75:6]};
  assign gzdLLzicase14914R2 = {gzdLLzilambda15508[139:70], gzdLLzilambda15508[145:140]};
  zdLLzicase14914  zdLLzicase14914R2 (gzdLLzicase14914R2[75:68], gzdLLzicase14914R2[67:60], gzdLLzicase14914R2[59:52], gzdLLzicase14914R2[51:44], gzdLLzicase14914R2[43:38], gzdLLzicase14914R2[37:21], gzdLLzicase14914R2[20:6], gzdLLzicase14914R2[5:0], callResR53);
  assign gzdLLzicase17968R8 = callResR53;
  zdLLzicase17968  zdLLzicase17968R8 (gzdLLzicase17968R8[69:0], callResR54);
  assign gzdLLzilambda19011 = callResR54;
  assign gzdLLzicase19009 = gzdLLzilambda19011[143:0];
  assign gzdLLzilambda15589 = gzdLLzicase19009[69:0];
  assign gzdLLzilambda19006 = {gzdLLzilambda15589[69:0], gzdLLzilambda15589[69:0]};
  assign gzdLLzicase18021R13 = gzdLLzilambda19006[139:0];
  zdLLzicase18021  zdLLzicase18021R13 (gzdLLzicase18021R13[139:70], gzdLLzicase18021R13[69:0], callResR55);
  assign gzdLLzilambda19001 = callResR55;
  assign gzdLLzicase18999 = gzdLLzilambda19001[143:0];
  assign gzdLLzilambda15587 = {gzdLLzicase18999[139:70], gzdLLzicase18999[69:0]};
  assign gMainzipcR3 = gzdLLzilambda15587[139:70];
  Mainzipc  MainzipcR3 (gMainzipcR3[69:0], callResR56);
  assign gzdLLzilambda18996 = {{7'h44{1'h0}}, callResR56, gzdLLzilambda15587[69:0]};
  assign gzdLLzicase18994 = gzdLLzilambda18996[143:0];
  assign gzdLLzilambda15585 = {gzdLLzicase18994[75:70], gzdLLzicase18994[69:0]};
  assign gzdLLzilambda15537 = {gzdLLzilambda15585[75:70], gzdLLzilambda15585[69:0]};
  assign gzdLLzilambda18917 = {gzdLLzilambda15537[69:0], gzdLLzilambda15537[69:0]};
  assign gzdLLzicase18021R14 = gzdLLzilambda18917[139:0];
  zdLLzicase18021  zdLLzicase18021R14 (gzdLLzicase18021R14[139:70], gzdLLzicase18021R14[69:0], callResR57);
  assign gzdLLzilambda18912 = {gzdLLzilambda15537[75:70], callResR57};
  assign gzdLLzicase18909 = {gzdLLzilambda18912[143:0], gzdLLzilambda18912[149:144]};
  assign gzdLLzilambda15535 = {gzdLLzicase18909[5:0], gzdLLzicase18909[145:76], gzdLLzicase18909[75:6]};
  assign gMainzioutputsR3 = gzdLLzilambda15535[139:70];
  Mainzioutputs  MainzioutputsR3 (gMainzioutputsR3[69:0], callResR58);
  assign gzdLLzilambda18905 = {gzdLLzilambda15535[145:140], {4'h5, {6'h37{1'h0}}}, callResR58, gzdLLzilambda15535[69:0]};
  assign gzdLLzicase18902 = {gzdLLzilambda18905[143:0], gzdLLzilambda18905[149:144]};
  assign gzdLLzilambda15532 = {gzdLLzicase18902[5:0], gzdLLzicase18902[90:76], gzdLLzicase18902[75:6]};
  assign gzdLLzicase14938R1 = {gzdLLzilambda15532[84:70], gzdLLzilambda15532[90:85]};
  zdLLzicase14938  zdLLzicase14938R1 (gzdLLzicase14938R1[20], gzdLLzicase14938R1[19:14], gzdLLzicase14938R1[13:6], gzdLLzicase14938R1[5:0], callResR59);
  assign gzdLLzilambda15524 = {callResR59, gzdLLzilambda15532[69:0]};
  assign gzdLLzilambda18898 = {gzdLLzilambda15524[69:0], gzdLLzilambda15524[69:0]};
  assign gzdLLzicase18021R15 = gzdLLzilambda18898[139:0];
  zdLLzicase18021  zdLLzicase18021R15 (gzdLLzicase18021R15[139:70], gzdLLzicase18021R15[69:0], callResR60);
  assign gzdLLzilambda18893 = {gzdLLzilambda15524[84:70], callResR60};
  assign gzdLLzicase18890 = {gzdLLzilambda18893[143:0], gzdLLzilambda18893[158:144]};
  assign gzdLLzilambda15522 = {gzdLLzicase18890[14:0], gzdLLzicase18890[154:85], gzdLLzicase18890[84:15]};
  assign gzdLLzicase14928R2 = {gzdLLzilambda15522[139:70], gzdLLzilambda15522[154:140]};
  zdLLzicase14928  zdLLzicase14928R2 (gzdLLzicase14928R2[84:77], gzdLLzicase14928R2[76:69], gzdLLzicase14928R2[68:61], gzdLLzicase14928R2[60:53], gzdLLzicase14928R2[52:47], gzdLLzicase14928R2[46:30], gzdLLzicase14928R2[29:15], gzdLLzicase14928R2[14:0], callResR61);
  assign gzdLLzicase17968R9 = callResR61;
  zdLLzicase17968  zdLLzicase17968R9 (gzdLLzicase17968R9[69:0], callResR62);
  assign gzdLLzilambda18991 = callResR62;
  assign gzdLLzicase18989 = gzdLLzilambda18991[143:0];
  assign gzdLLzilambda15583 = gzdLLzicase18989[69:0];
  assign gzdLLzilambda18986 = {gzdLLzilambda15583[69:0], gzdLLzilambda15583[69:0]};
  assign gzdLLzicase18021R16 = gzdLLzilambda18986[139:0];
  zdLLzicase18021  zdLLzicase18021R16 (gzdLLzicase18021R16[139:70], gzdLLzicase18021R16[69:0], callResR63);
  assign gzdLLzilambda18981 = callResR63;
  assign gzdLLzicase18979 = gzdLLzilambda18981[143:0];
  assign gzdLLzilambda15581 = {gzdLLzicase18979[139:70], gzdLLzicase18979[69:0]};
  assign gMainzioutputsR4 = gzdLLzilambda15581[139:70];
  Mainzioutputs  MainzioutputsR4 (gMainzioutputsR4[69:0], callResR64);
  assign gzdLLzilambda18976 = {{4'h5, {6'h37{1'h0}}}, callResR64, gzdLLzilambda15581[69:0]};
  assign gzdLLzicase18974 = gzdLLzilambda18976[143:0];
  assign gzdLLzilambda15579 = {gzdLLzicase18974[84:70], gzdLLzicase18974[69:0]};
  assign gzdLLzicase14964R1 = gzdLLzilambda15579[84:70];
  zdLLzicase14964  zdLLzicase14964R1 (gzdLLzicase14964R1[14], gzdLLzicase14964R1[13:8], gzdLLzicase14964R1[7:0], callResR65);
  assign gzdLLzilambda15551 = {callResR65, gzdLLzilambda15579[69:0]};
  assign gzdLLzilambda18934 = {gzdLLzilambda15551[69:0], gzdLLzilambda15551[69:0]};
  assign gzdLLzicase18021R17 = gzdLLzilambda18934[139:0];
  zdLLzicase18021  zdLLzicase18021R17 (gzdLLzicase18021R17[139:70], gzdLLzicase18021R17[69:0], callResR66);
  assign gzdLLzilambda18929 = {gzdLLzilambda15551[84:70], callResR66};
  assign gzdLLzicase18926 = {gzdLLzilambda18929[143:0], gzdLLzilambda18929[158:144]};
  assign gzdLLzilambda15549 = {gzdLLzicase18926[14:0], gzdLLzicase18926[154:85], gzdLLzicase18926[84:15]};
  assign gzdLLzicase14928R3 = {gzdLLzilambda15549[139:70], gzdLLzilambda15549[154:140]};
  zdLLzicase14928  zdLLzicase14928R3 (gzdLLzicase14928R3[84:77], gzdLLzicase14928R3[76:69], gzdLLzicase14928R3[68:61], gzdLLzicase14928R3[60:53], gzdLLzicase14928R3[52:47], gzdLLzicase14928R3[46:30], gzdLLzicase14928R3[29:15], gzdLLzicase14928R3[14:0], callResR67);
  assign gzdLLzicase17968R10 = callResR67;
  zdLLzicase17968  zdLLzicase17968R10 (gzdLLzicase17968R10[69:0], callResR68);
  assign gzdLLzilambda18971 = callResR68;
  assign gzdLLzicase18969 = gzdLLzilambda18971[143:0];
  assign gzdLLzilambda15577 = gzdLLzicase18969[69:0];
  assign gzdLLzilambda18966 = {gzdLLzilambda15577[69:0], gzdLLzilambda15577[69:0]};
  assign gzdLLzicase18021R18 = gzdLLzilambda18966[139:0];
  zdLLzicase18021  zdLLzicase18021R18 (gzdLLzicase18021R18[139:70], gzdLLzicase18021R18[69:0], callResR69);
  assign gzdLLzilambda18961 = callResR69;
  assign gzdLLzicase18959 = gzdLLzilambda18961[143:0];
  assign gzdLLzilambda15575 = {gzdLLzicase18959[139:70], gzdLLzicase18959[69:0]};
  assign gMainzioutputsR5 = gzdLLzilambda15575[139:70];
  Mainzioutputs  MainzioutputsR5 (gMainzioutputsR5[69:0], callResR70);
  assign gzdLLzilambda18956 = {{4'h5, {6'h37{1'h0}}}, callResR70, gzdLLzilambda15575[69:0]};
  assign gzdLLzicase18954 = gzdLLzilambda18956[143:0];
  assign gzdLLzilambda15573 = {gzdLLzicase18954[84:70], gzdLLzicase18954[69:0]};
  assign gzdLLzicase15741 = {gzdLLzilambda15749[148:140], gzdLLzilambda15749[69:0]};
  assign gzdLLzilambda15407 = {gzdLLzicase15741[75:70], gzdLLzicase15741[69:0]};
  assign gzdLLzilambda18836 = {gzdLLzilambda15407[69:0], gzdLLzilambda15407[69:0]};
  assign gzdLLzilambda15200R3 = gzdLLzilambda18836[139:0];
  zdLLzilambda15200  zdLLzilambda15200R3 (gzdLLzilambda15200R3[139:70], gzdLLzilambda15200R3[69:0], callResR71);
  assign gzdLLzilambda18831 = callResR71;
  assign gzdLLzicase17888R9 = gzdLLzilambda18831[77:0];
  zdLLzicase17888  zdLLzicase17888R9 (gzdLLzicase17888R9[77:70], gzdLLzicase17888R9[69:0], callResR72);
  assign gzdLLzilambda18826 = {gzdLLzilambda15407[75:70], callResR72};
  assign gzdLLzicase18823 = {gzdLLzilambda18826[143:0], gzdLLzilambda18826[149:144]};
  assign gzdLLzilambda15405 = {gzdLLzicase18823[5:0], gzdLLzicase18823[83:76], gzdLLzicase18823[75:6]};
  assign gzdLLzilambda15227 = {gzdLLzilambda15405[83:78], gzdLLzilambda15405[69:0]};
  assign gzdLLzilambda18535 = {gzdLLzilambda15227[69:0], gzdLLzilambda15227[69:0]};
  assign gzdLLzicase18021R19 = gzdLLzilambda18535[139:0];
  zdLLzicase18021  zdLLzicase18021R19 (gzdLLzicase18021R19[139:70], gzdLLzicase18021R19[69:0], callResR73);
  assign gzdLLzilambda18530 = {gzdLLzilambda15227[75:70], callResR73};
  assign gzdLLzicase18527 = {gzdLLzilambda18530[143:0], gzdLLzilambda18530[149:144]};
  assign gzdLLzilambda15225 = {gzdLLzicase18527[5:0], gzdLLzicase18527[145:76], gzdLLzicase18527[75:6]};
  assign gMainzioutputsR6 = gzdLLzilambda15225[139:70];
  Mainzioutputs  MainzioutputsR6 (gMainzioutputsR6[69:0], callResR74);
  assign gzdLLzilambda18523 = {gzdLLzilambda15225[145:140], {4'h5, {6'h37{1'h0}}}, callResR74, gzdLLzilambda15225[69:0]};
  assign gzdLLzicase18520 = {gzdLLzilambda18523[143:0], gzdLLzilambda18523[149:144]};
  assign gzdLLzilambda15222 = {gzdLLzicase18520[5:0], gzdLLzicase18520[90:76], gzdLLzicase18520[75:6]};
  assign gzdLLzicase14938R2 = {gzdLLzilambda15222[84:70], gzdLLzilambda15222[90:85]};
  zdLLzicase14938  zdLLzicase14938R2 (gzdLLzicase14938R2[20], gzdLLzicase14938R2[19:14], gzdLLzicase14938R2[13:6], gzdLLzicase14938R2[5:0], callResR75);
  assign gzdLLzilambda15214 = {callResR75, gzdLLzilambda15222[69:0]};
  assign gzdLLzilambda18516 = {gzdLLzilambda15214[69:0], gzdLLzilambda15214[69:0]};
  assign gzdLLzicase18021R20 = gzdLLzilambda18516[139:0];
  zdLLzicase18021  zdLLzicase18021R20 (gzdLLzicase18021R20[139:70], gzdLLzicase18021R20[69:0], callResR76);
  assign gzdLLzilambda18511 = {gzdLLzilambda15214[84:70], callResR76};
  assign gzdLLzicase18508 = {gzdLLzilambda18511[143:0], gzdLLzilambda18511[158:144]};
  assign gzdLLzilambda15212 = {gzdLLzicase18508[14:0], gzdLLzicase18508[154:85], gzdLLzicase18508[84:15]};
  assign gzdLLzicase14928R4 = {gzdLLzilambda15212[139:70], gzdLLzilambda15212[154:140]};
  zdLLzicase14928  zdLLzicase14928R4 (gzdLLzicase14928R4[84:77], gzdLLzicase14928R4[76:69], gzdLLzicase14928R4[68:61], gzdLLzicase14928R4[60:53], gzdLLzicase14928R4[52:47], gzdLLzicase14928R4[46:30], gzdLLzicase14928R4[29:15], gzdLLzicase14928R4[14:0], callResR77);
  assign gzdLLzicase17968R11 = callResR77;
  zdLLzicase17968  zdLLzicase17968R11 (gzdLLzicase17968R11[69:0], callResR78);
  assign gzdLLzilambda18819 = {gzdLLzilambda15405[77:70], callResR78};
  assign gzdLLzicase18816 = {gzdLLzilambda18819[143:0], gzdLLzilambda18819[151:144]};
  assign gzdLLzilambda15402 = {gzdLLzicase18816[7:0], gzdLLzicase18816[77:8]};
  assign gzdLLzilambda15254 = {gzdLLzilambda15402[77:70], gzdLLzilambda15402[69:0]};
  assign gzdLLzilambda18571 = {gzdLLzilambda15254[69:0], gzdLLzilambda15254[69:0]};
  assign gzdLLzicase18021R21 = gzdLLzilambda18571[139:0];
  zdLLzicase18021  zdLLzicase18021R21 (gzdLLzicase18021R21[139:70], gzdLLzicase18021R21[69:0], callResR79);
  assign gzdLLzilambda18566 = {gzdLLzilambda15254[77:70], callResR79};
  assign gzdLLzicase18563 = {gzdLLzilambda18566[143:0], gzdLLzilambda18566[151:144]};
  assign gzdLLzilambda15252 = {gzdLLzicase18563[7:0], gzdLLzicase18563[147:78], gzdLLzicase18563[77:8]};
  assign gMainzioutputsR7 = gzdLLzilambda15252[139:70];
  Mainzioutputs  MainzioutputsR7 (gMainzioutputsR7[69:0], callResR80);
  assign gzdLLzilambda18559 = {gzdLLzilambda15252[147:140], {4'h5, {6'h37{1'h0}}}, callResR80, gzdLLzilambda15252[69:0]};
  assign gzdLLzicase18556 = {gzdLLzilambda18559[143:0], gzdLLzilambda18559[151:144]};
  assign gzdLLzilambda15249 = {gzdLLzicase18556[7:0], gzdLLzicase18556[92:78], gzdLLzicase18556[77:8]};
  assign gzdLLzicase15246 = {gzdLLzilambda15249[84:70], gzdLLzilambda15249[92:85]};
  assign gzdLLzilambda15241 = {{gzdLLzicase15246[22], gzdLLzicase15246[21:16], gzdLLzicase15246[7:0]}, gzdLLzilambda15249[69:0]};
  assign gzdLLzilambda18552 = {gzdLLzilambda15241[69:0], gzdLLzilambda15241[69:0]};
  assign gzdLLzicase18021R22 = gzdLLzilambda18552[139:0];
  zdLLzicase18021  zdLLzicase18021R22 (gzdLLzicase18021R22[139:70], gzdLLzicase18021R22[69:0], callResR81);
  assign gzdLLzilambda18547 = {gzdLLzilambda15241[84:70], callResR81};
  assign gzdLLzicase18544 = {gzdLLzilambda18547[143:0], gzdLLzilambda18547[158:144]};
  assign gzdLLzilambda15239 = {gzdLLzicase18544[14:0], gzdLLzicase18544[154:85], gzdLLzicase18544[84:15]};
  assign gzdLLzicase14928R5 = {gzdLLzilambda15239[139:70], gzdLLzilambda15239[154:140]};
  zdLLzicase14928  zdLLzicase14928R5 (gzdLLzicase14928R5[84:77], gzdLLzicase14928R5[76:69], gzdLLzicase14928R5[68:61], gzdLLzicase14928R5[60:53], gzdLLzicase14928R5[52:47], gzdLLzicase14928R5[46:30], gzdLLzicase14928R5[29:15], gzdLLzicase14928R5[14:0], callResR82);
  assign gzdLLzicase17968R12 = callResR82;
  zdLLzicase17968  zdLLzicase17968R12 (gzdLLzicase17968R12[69:0], callResR83);
  assign gzdLLzilambda18812 = callResR83;
  assign gzdLLzicase18810 = gzdLLzilambda18812[143:0];
  assign gzdLLzilambda15399 = gzdLLzicase18810[69:0];
  assign gzdLLzilambda18807 = {gzdLLzilambda15399[69:0], gzdLLzilambda15399[69:0]};
  assign gzdLLzicase18021R23 = gzdLLzilambda18807[139:0];
  zdLLzicase18021  zdLLzicase18021R23 (gzdLLzicase18021R23[139:70], gzdLLzicase18021R23[69:0], callResR84);
  assign gzdLLzilambda18802 = callResR84;
  assign gzdLLzicase18800 = gzdLLzilambda18802[143:0];
  assign gzdLLzilambda15397 = {gzdLLzicase18800[139:70], gzdLLzicase18800[69:0]};
  assign gMainzioutputsR8 = gzdLLzilambda15397[139:70];
  Mainzioutputs  MainzioutputsR8 (gMainzioutputsR8[69:0], callResR85);
  assign gzdLLzilambda18797 = {{4'h5, {6'h37{1'h0}}}, callResR85, gzdLLzilambda15397[69:0]};
  assign gzdLLzicase18795 = gzdLLzilambda18797[143:0];
  assign gzdLLzilambda15395 = {gzdLLzicase18795[84:70], gzdLLzicase18795[69:0]};
  assign gzdLLzicase15272 = gzdLLzilambda15395[84:70];
  assign gzdLLzilambda15268 = {{1'h1, gzdLLzicase15272[13:8], gzdLLzicase15272[7:0]}, gzdLLzilambda15395[69:0]};
  assign gzdLLzilambda18588 = {gzdLLzilambda15268[69:0], gzdLLzilambda15268[69:0]};
  assign gzdLLzicase18021R24 = gzdLLzilambda18588[139:0];
  zdLLzicase18021  zdLLzicase18021R24 (gzdLLzicase18021R24[139:70], gzdLLzicase18021R24[69:0], callResR86);
  assign gzdLLzilambda18583 = {gzdLLzilambda15268[84:70], callResR86};
  assign gzdLLzicase18580 = {gzdLLzilambda18583[143:0], gzdLLzilambda18583[158:144]};
  assign gzdLLzilambda15266 = {gzdLLzicase18580[14:0], gzdLLzicase18580[154:85], gzdLLzicase18580[84:15]};
  assign gzdLLzicase14928R6 = {gzdLLzilambda15266[139:70], gzdLLzilambda15266[154:140]};
  zdLLzicase14928  zdLLzicase14928R6 (gzdLLzicase14928R6[84:77], gzdLLzicase14928R6[76:69], gzdLLzicase14928R6[68:61], gzdLLzicase14928R6[60:53], gzdLLzicase14928R6[52:47], gzdLLzicase14928R6[46:30], gzdLLzicase14928R6[29:15], gzdLLzicase14928R6[14:0], callResR87);
  assign gzdLLzicase17968R13 = callResR87;
  zdLLzicase17968  zdLLzicase17968R13 (gzdLLzicase17968R13[69:0], callResR88);
  assign gzdLLzilambda18792 = callResR88;
  assign gzdLLzicase18790 = gzdLLzilambda18792[143:0];
  assign gzdLLzilambda15393 = gzdLLzicase18790[69:0];
  assign gzdLLzilambda18787 = {gzdLLzilambda15393[69:0], gzdLLzilambda15393[69:0]};
  assign gzdLLzicase18021R25 = gzdLLzilambda18787[139:0];
  zdLLzicase18021  zdLLzicase18021R25 (gzdLLzicase18021R25[139:70], gzdLLzicase18021R25[69:0], callResR89);
  assign gzdLLzilambda18782 = callResR89;
  assign gzdLLzicase18780 = gzdLLzilambda18782[143:0];
  assign gzdLLzilambda15391 = {gzdLLzicase18780[139:70], gzdLLzicase18780[69:0]};
  assign gMainzioutputsR9 = gzdLLzilambda15391[139:70];
  Mainzioutputs  MainzioutputsR9 (gMainzioutputsR9[69:0], callResR90);
  assign gzdLLzilambda18777 = {{4'h5, {6'h37{1'h0}}}, callResR90, gzdLLzilambda15391[69:0]};
  assign gzdLLzicase18775 = gzdLLzilambda18777[143:0];
  assign gzdLLzilambda15389 = {gzdLLzicase18775[84:70], gzdLLzicase18775[69:0]};
  assign gzdLLzicase15743 = {gzdLLzilambda15749[148:140], gzdLLzilambda15749[69:0]};
  assign gzdLLzilambda15198 = {gzdLLzicase15743[75:70], gzdLLzicase15743[69:0]};
  assign gzdLLzilambda15029 = {gzdLLzilambda15198[75:70], gzdLLzilambda15198[69:0]};
  assign gzdLLzilambda18221 = {gzdLLzilambda15029[69:0], gzdLLzilambda15029[69:0]};
  assign gzdLLzicase18021R26 = gzdLLzilambda18221[139:0];
  zdLLzicase18021  zdLLzicase18021R26 (gzdLLzicase18021R26[139:70], gzdLLzicase18021R26[69:0], callResR91);
  assign gzdLLzilambda18216 = {gzdLLzilambda15029[75:70], callResR91};
  assign gzdLLzicase18213 = {gzdLLzilambda18216[143:0], gzdLLzilambda18216[149:144]};
  assign gzdLLzilambda15027 = {gzdLLzicase18213[5:0], gzdLLzicase18213[145:76], gzdLLzicase18213[75:6]};
  assign gMainzioutputsR10 = gzdLLzilambda15027[139:70];
  Mainzioutputs  MainzioutputsR10 (gMainzioutputsR10[69:0], callResR92);
  assign gzdLLzilambda18209 = {gzdLLzilambda15027[145:140], {4'h5, {6'h37{1'h0}}}, callResR92, gzdLLzilambda15027[69:0]};
  assign gzdLLzicase18206 = {gzdLLzilambda18209[143:0], gzdLLzilambda18209[149:144]};
  assign gzdLLzilambda15024 = {gzdLLzicase18206[5:0], gzdLLzicase18206[90:76], gzdLLzicase18206[75:6]};
  assign gzdLLzicase14938R3 = {gzdLLzilambda15024[84:70], gzdLLzilambda15024[90:85]};
  zdLLzicase14938  zdLLzicase14938R3 (gzdLLzicase14938R3[20], gzdLLzicase14938R3[19:14], gzdLLzicase14938R3[13:6], gzdLLzicase14938R3[5:0], callResR93);
  assign gzdLLzilambda15016 = {callResR93, gzdLLzilambda15024[69:0]};
  assign gzdLLzilambda18202 = {gzdLLzilambda15016[69:0], gzdLLzilambda15016[69:0]};
  assign gzdLLzicase18021R27 = gzdLLzilambda18202[139:0];
  zdLLzicase18021  zdLLzicase18021R27 (gzdLLzicase18021R27[139:70], gzdLLzicase18021R27[69:0], callResR94);
  assign gzdLLzilambda18197 = {gzdLLzilambda15016[84:70], callResR94};
  assign gzdLLzicase18194 = {gzdLLzilambda18197[143:0], gzdLLzilambda18197[158:144]};
  assign gzdLLzilambda15014 = {gzdLLzicase18194[14:0], gzdLLzicase18194[154:85], gzdLLzicase18194[84:15]};
  assign gzdLLzicase14928R7 = {gzdLLzilambda15014[139:70], gzdLLzilambda15014[154:140]};
  zdLLzicase14928  zdLLzicase14928R7 (gzdLLzicase14928R7[84:77], gzdLLzicase14928R7[76:69], gzdLLzicase14928R7[68:61], gzdLLzicase14928R7[60:53], gzdLLzicase14928R7[52:47], gzdLLzicase14928R7[46:30], gzdLLzicase14928R7[29:15], gzdLLzicase14928R7[14:0], callResR95);
  assign gzdLLzicase17968R14 = callResR95;
  zdLLzicase17968  zdLLzicase17968R14 (gzdLLzicase17968R14[69:0], callResR96);
  assign gzdLLzilambda18499 = callResR96;
  assign gzdLLzicase18497 = gzdLLzilambda18499[143:0];
  assign gzdLLzilambda15196 = gzdLLzicase18497[69:0];
  assign gzdLLzilambda18494 = {gzdLLzilambda15196[69:0], gzdLLzilambda15196[69:0]};
  assign gzdLLzicase18021R28 = gzdLLzilambda18494[139:0];
  zdLLzicase18021  zdLLzicase18021R28 (gzdLLzicase18021R28[139:70], gzdLLzicase18021R28[69:0], callResR97);
  assign gzdLLzilambda18489 = callResR97;
  assign gzdLLzicase18487 = gzdLLzilambda18489[143:0];
  assign gzdLLzilambda15194 = {gzdLLzicase18487[139:70], gzdLLzicase18487[69:0]};
  assign gMainzioutputsR11 = gzdLLzilambda15194[139:70];
  Mainzioutputs  MainzioutputsR11 (gMainzioutputsR11[69:0], callResR98);
  assign gzdLLzilambda18484 = {{4'h5, {6'h37{1'h0}}}, callResR98, gzdLLzilambda15194[69:0]};
  assign gzdLLzicase18482 = gzdLLzilambda18484[143:0];
  assign gzdLLzilambda15192 = {gzdLLzicase18482[84:70], gzdLLzicase18482[69:0]};
  assign gzdLLzicase14964R2 = gzdLLzilambda15192[84:70];
  zdLLzicase14964  zdLLzicase14964R2 (gzdLLzicase14964R2[14], gzdLLzicase14964R2[13:8], gzdLLzicase14964R2[7:0], callResR99);
  assign gzdLLzilambda15043 = {callResR99, gzdLLzilambda15192[69:0]};
  assign gzdLLzilambda18238 = {gzdLLzilambda15043[69:0], gzdLLzilambda15043[69:0]};
  assign gzdLLzicase18021R29 = gzdLLzilambda18238[139:0];
  zdLLzicase18021  zdLLzicase18021R29 (gzdLLzicase18021R29[139:70], gzdLLzicase18021R29[69:0], callResR100);
  assign gzdLLzilambda18233 = {gzdLLzilambda15043[84:70], callResR100};
  assign gzdLLzicase18230 = {gzdLLzilambda18233[143:0], gzdLLzilambda18233[158:144]};
  assign gzdLLzilambda15041 = {gzdLLzicase18230[14:0], gzdLLzicase18230[154:85], gzdLLzicase18230[84:15]};
  assign gzdLLzicase14928R8 = {gzdLLzilambda15041[139:70], gzdLLzilambda15041[154:140]};
  zdLLzicase14928  zdLLzicase14928R8 (gzdLLzicase14928R8[84:77], gzdLLzicase14928R8[76:69], gzdLLzicase14928R8[68:61], gzdLLzicase14928R8[60:53], gzdLLzicase14928R8[52:47], gzdLLzicase14928R8[46:30], gzdLLzicase14928R8[29:15], gzdLLzicase14928R8[14:0], callResR101);
  assign gzdLLzicase17968R15 = callResR101;
  zdLLzicase17968  zdLLzicase17968R15 (gzdLLzicase17968R15[69:0], callResR102);
  assign gzdLLzilambda18479 = callResR102;
  assign gzdLLzicase18477 = gzdLLzilambda18479[143:0];
  assign gzdLLzilambda15190 = gzdLLzicase18477[69:0];
  assign gzdLLzilambda18474 = {gzdLLzilambda15190[69:0], gzdLLzilambda15190[69:0]};
  assign gzdLLzicase18021R30 = gzdLLzilambda18474[139:0];
  zdLLzicase18021  zdLLzicase18021R30 (gzdLLzicase18021R30[139:70], gzdLLzicase18021R30[69:0], callResR103);
  assign gzdLLzilambda18469 = callResR103;
  assign gzdLLzicase18467 = gzdLLzilambda18469[143:0];
  assign gzdLLzilambda15188 = {gzdLLzicase18467[139:70], gzdLLzicase18467[69:0]};
  assign gMainzioutputsR12 = gzdLLzilambda15188[139:70];
  Mainzioutputs  MainzioutputsR12 (gMainzioutputsR12[69:0], callResR104);
  assign gzdLLzilambda18464 = {{4'h5, {6'h37{1'h0}}}, callResR104, gzdLLzilambda15188[69:0]};
  assign gzdLLzicase18462 = gzdLLzilambda18464[143:0];
  assign gzdLLzilambda15186 = {gzdLLzicase18462[84:70], gzdLLzicase18462[69:0]};
  assign gzdLLzicase19261 = {gzdLLzilambda15749[148:140], gzdLLzilambda15749[69:0]};
  assign gzdLLzicase15744 = gzdLLzicase19261[69:0];
  assign gzdLLzilambda18033 = {gzdLLzicase15744[69:0], gzdLLzicase15744[69:0]};
  assign gzdLLzicase18021R31 = gzdLLzilambda18033[139:0];
  zdLLzicase18021  zdLLzicase18021R31 (gzdLLzicase18021R31[139:70], gzdLLzicase18021R31[69:0], callResR105);
  assign gzdLLzilambda18028 = callResR105;
  assign gzdLLzicase18026 = gzdLLzilambda18028[143:0];
  assign gzdLLzilambda15002 = {gzdLLzicase18026[139:70], gzdLLzicase18026[69:0]};
  assign gMainzipcR4 = gzdLLzilambda15002[139:70];
  Mainzipc  MainzipcR4 (gMainzipcR4[69:0], callResR106);
  assign gzdLLzilambda18185 = {{7'h44{1'h0}}, callResR106, gzdLLzilambda15002[69:0]};
  assign gzdLLzicase18183 = gzdLLzilambda18185[143:0];
  assign gzdLLzilambda15000 = {gzdLLzicase18183[75:70], gzdLLzicase18183[69:0]};
  assign binOpR5 = {gzdLLzilambda15000[75:70], 6'h01};
  assign gzdLLzilambda14919 = {binOpR5[11:6] + binOpR5[5:0], gzdLLzilambda15000[69:0]};
  assign gzdLLzilambda18050 = {gzdLLzilambda14919[69:0], gzdLLzilambda14919[69:0]};
  assign gzdLLzicase18021R32 = gzdLLzilambda18050[139:0];
  zdLLzicase18021  zdLLzicase18021R32 (gzdLLzicase18021R32[139:70], gzdLLzicase18021R32[69:0], callResR107);
  assign gzdLLzilambda18045 = {gzdLLzilambda14919[75:70], callResR107};
  assign gzdLLzicase18042 = {gzdLLzilambda18045[143:0], gzdLLzilambda18045[149:144]};
  assign gzdLLzilambda14917 = {gzdLLzicase18042[5:0], gzdLLzicase18042[145:76], gzdLLzicase18042[75:6]};
  assign gzdLLzicase14914R3 = {gzdLLzilambda14917[139:70], gzdLLzilambda14917[145:140]};
  zdLLzicase14914  zdLLzicase14914R3 (gzdLLzicase14914R3[75:68], gzdLLzicase14914R3[67:60], gzdLLzicase14914R3[59:52], gzdLLzicase14914R3[51:44], gzdLLzicase14914R3[43:38], gzdLLzicase14914R3[37:21], gzdLLzicase14914R3[20:6], gzdLLzicase14914R3[5:0], callResR108);
  assign gzdLLzicase17968R16 = callResR108;
  zdLLzicase17968  zdLLzicase17968R16 (gzdLLzicase17968R16[69:0], callResR109);
  assign gzdLLzilambda18180 = callResR109;
  assign gzdLLzicase18178 = gzdLLzilambda18180[143:0];
  assign gzdLLzilambda14998 = gzdLLzicase18178[69:0];
  assign gzdLLzilambda18175 = {gzdLLzilambda14998[69:0], gzdLLzilambda14998[69:0]};
  assign gzdLLzicase18021R33 = gzdLLzilambda18175[139:0];
  zdLLzicase18021  zdLLzicase18021R33 (gzdLLzicase18021R33[139:70], gzdLLzicase18021R33[69:0], callResR110);
  assign gzdLLzilambda18170 = callResR110;
  assign gzdLLzicase18168 = gzdLLzilambda18170[143:0];
  assign gzdLLzilambda14996 = {gzdLLzicase18168[139:70], gzdLLzicase18168[69:0]};
  assign gMainzipcR5 = gzdLLzilambda14996[139:70];
  Mainzipc  MainzipcR5 (gMainzipcR5[69:0], callResR111);
  assign gzdLLzilambda18165 = {{7'h44{1'h0}}, callResR111, gzdLLzilambda14996[69:0]};
  assign gzdLLzicase18163 = gzdLLzilambda18165[143:0];
  assign gzdLLzilambda14994 = {gzdLLzicase18163[75:70], gzdLLzicase18163[69:0]};
  assign gzdLLzilambda14946 = {gzdLLzilambda14994[75:70], gzdLLzilambda14994[69:0]};
  assign gzdLLzilambda18086 = {gzdLLzilambda14946[69:0], gzdLLzilambda14946[69:0]};
  assign gzdLLzicase18021R34 = gzdLLzilambda18086[139:0];
  zdLLzicase18021  zdLLzicase18021R34 (gzdLLzicase18021R34[139:70], gzdLLzicase18021R34[69:0], callResR112);
  assign gzdLLzilambda18081 = {gzdLLzilambda14946[75:70], callResR112};
  assign gzdLLzicase18078 = {gzdLLzilambda18081[143:0], gzdLLzilambda18081[149:144]};
  assign gzdLLzilambda14944 = {gzdLLzicase18078[5:0], gzdLLzicase18078[145:76], gzdLLzicase18078[75:6]};
  assign gMainzioutputsR13 = gzdLLzilambda14944[139:70];
  Mainzioutputs  MainzioutputsR13 (gMainzioutputsR13[69:0], callResR113);
  assign gzdLLzilambda18074 = {gzdLLzilambda14944[145:140], {4'h5, {6'h37{1'h0}}}, callResR113, gzdLLzilambda14944[69:0]};
  assign gzdLLzicase18071 = {gzdLLzilambda18074[143:0], gzdLLzilambda18074[149:144]};
  assign gzdLLzilambda14941 = {gzdLLzicase18071[5:0], gzdLLzicase18071[90:76], gzdLLzicase18071[75:6]};
  assign gzdLLzicase14938R4 = {gzdLLzilambda14941[84:70], gzdLLzilambda14941[90:85]};
  zdLLzicase14938  zdLLzicase14938R4 (gzdLLzicase14938R4[20], gzdLLzicase14938R4[19:14], gzdLLzicase14938R4[13:6], gzdLLzicase14938R4[5:0], callResR114);
  assign gzdLLzilambda14933 = {callResR114, gzdLLzilambda14941[69:0]};
  assign gzdLLzilambda18067 = {gzdLLzilambda14933[69:0], gzdLLzilambda14933[69:0]};
  assign gzdLLzicase18021R35 = gzdLLzilambda18067[139:0];
  zdLLzicase18021  zdLLzicase18021R35 (gzdLLzicase18021R35[139:70], gzdLLzicase18021R35[69:0], callResR115);
  assign gzdLLzilambda18062 = {gzdLLzilambda14933[84:70], callResR115};
  assign gzdLLzicase18059 = {gzdLLzilambda18062[143:0], gzdLLzilambda18062[158:144]};
  assign gzdLLzilambda14931 = {gzdLLzicase18059[14:0], gzdLLzicase18059[154:85], gzdLLzicase18059[84:15]};
  assign gzdLLzicase14928R9 = {gzdLLzilambda14931[139:70], gzdLLzilambda14931[154:140]};
  zdLLzicase14928  zdLLzicase14928R9 (gzdLLzicase14928R9[84:77], gzdLLzicase14928R9[76:69], gzdLLzicase14928R9[68:61], gzdLLzicase14928R9[60:53], gzdLLzicase14928R9[52:47], gzdLLzicase14928R9[46:30], gzdLLzicase14928R9[29:15], gzdLLzicase14928R9[14:0], callResR116);
  assign gzdLLzicase17968R17 = callResR116;
  zdLLzicase17968  zdLLzicase17968R17 (gzdLLzicase17968R17[69:0], callResR117);
  assign gzdLLzilambda18160 = callResR117;
  assign gzdLLzicase18158 = gzdLLzilambda18160[143:0];
  assign gzdLLzilambda14992 = gzdLLzicase18158[69:0];
  assign gzdLLzilambda18155 = {gzdLLzilambda14992[69:0], gzdLLzilambda14992[69:0]};
  assign gzdLLzicase18021R36 = gzdLLzilambda18155[139:0];
  zdLLzicase18021  zdLLzicase18021R36 (gzdLLzicase18021R36[139:70], gzdLLzicase18021R36[69:0], callResR118);
  assign gzdLLzilambda18150 = callResR118;
  assign gzdLLzicase18148 = gzdLLzilambda18150[143:0];
  assign gzdLLzilambda14990 = {gzdLLzicase18148[139:70], gzdLLzicase18148[69:0]};
  assign gMainzioutputsR14 = gzdLLzilambda14990[139:70];
  Mainzioutputs  MainzioutputsR14 (gMainzioutputsR14[69:0], callResR119);
  assign gzdLLzilambda18145 = {{4'h5, {6'h37{1'h0}}}, callResR119, gzdLLzilambda14990[69:0]};
  assign gzdLLzicase18143 = gzdLLzilambda18145[143:0];
  assign gzdLLzilambda14988 = {gzdLLzicase18143[84:70], gzdLLzicase18143[69:0]};
  assign gzdLLzicase14964R3 = gzdLLzilambda14988[84:70];
  zdLLzicase14964  zdLLzicase14964R3 (gzdLLzicase14964R3[14], gzdLLzicase14964R3[13:8], gzdLLzicase14964R3[7:0], callResR120);
  assign gzdLLzilambda14960 = {callResR120, gzdLLzilambda14988[69:0]};
  assign gzdLLzilambda18103 = {gzdLLzilambda14960[69:0], gzdLLzilambda14960[69:0]};
  assign gzdLLzicase18021R37 = gzdLLzilambda18103[139:0];
  zdLLzicase18021  zdLLzicase18021R37 (gzdLLzicase18021R37[139:70], gzdLLzicase18021R37[69:0], callResR121);
  assign gzdLLzilambda18098 = {gzdLLzilambda14960[84:70], callResR121};
  assign gzdLLzicase18095 = {gzdLLzilambda18098[143:0], gzdLLzilambda18098[158:144]};
  assign gzdLLzilambda14958 = {gzdLLzicase18095[14:0], gzdLLzicase18095[154:85], gzdLLzicase18095[84:15]};
  assign gzdLLzicase14928R10 = {gzdLLzilambda14958[139:70], gzdLLzilambda14958[154:140]};
  zdLLzicase14928  zdLLzicase14928R10 (gzdLLzicase14928R10[84:77], gzdLLzicase14928R10[76:69], gzdLLzicase14928R10[68:61], gzdLLzicase14928R10[60:53], gzdLLzicase14928R10[52:47], gzdLLzicase14928R10[46:30], gzdLLzicase14928R10[29:15], gzdLLzicase14928R10[14:0], callResR122);
  assign gzdLLzicase17968R18 = callResR122;
  zdLLzicase17968  zdLLzicase17968R18 (gzdLLzicase17968R18[69:0], callResR123);
  assign gzdLLzilambda18140 = callResR123;
  assign gzdLLzicase18138 = gzdLLzilambda18140[143:0];
  assign gzdLLzilambda14986 = gzdLLzicase18138[69:0];
  assign gzdLLzilambda18135 = {gzdLLzilambda14986[69:0], gzdLLzilambda14986[69:0]};
  assign gzdLLzicase18021R38 = gzdLLzilambda18135[139:0];
  zdLLzicase18021  zdLLzicase18021R38 (gzdLLzicase18021R38[139:70], gzdLLzicase18021R38[69:0], callResR124);
  assign gzdLLzilambda18130 = callResR124;
  assign gzdLLzicase18128 = gzdLLzilambda18130[143:0];
  assign gzdLLzilambda14984 = {gzdLLzicase18128[139:70], gzdLLzicase18128[69:0]};
  assign gMainzioutputsR15 = gzdLLzilambda14984[139:70];
  Mainzioutputs  MainzioutputsR15 (gMainzioutputsR15[69:0], callResR125);
  assign gzdLLzilambda18125 = {{4'h5, {6'h37{1'h0}}}, callResR125, gzdLLzilambda14984[69:0]};
  assign gzdLLzicase18123 = gzdLLzilambda18125[143:0];
  assign gzdLLzilambda14982 = {gzdLLzicase18123[84:70], gzdLLzicase18123[69:0]};
  assign gzdLLzilambda19245 = (gzdLLzicase19261[78:76] == 3'h0) ? {{1'h1, {6'h36{1'h0}}}, gzdLLzilambda14982[84:70], 4'h0, gzdLLzilambda14982[69:0]} : ((gzdLLzicase15743[78:76] == 3'h1) ? {{1'h1, {6'h36{1'h0}}}, gzdLLzilambda15186[84:70], 4'h2, gzdLLzilambda15186[69:0]} : ((gzdLLzicase15741[78:76] == 3'h2) ? {{1'h1, {6'h36{1'h0}}}, gzdLLzilambda15389[84:70], 4'h4, gzdLLzilambda15389[69:0]} : ((gzdLLzicase15739[78:76] == 3'h3) ? {{1'h1, {6'h36{1'h0}}}, gzdLLzilambda15573[84:70], 4'h5, gzdLLzilambda15573[69:0]} : {{1'h1, {6'h36{1'h0}}}, gzdLLzilambda15712[84:70], 4'h6, gzdLLzilambda15712[69:0]})));
  assign gzdLLzicase19243 = gzdLLzilambda19245[143:0];
  zdLLzicase19243  zdLLzicase19243 (gzdLLzicase19243[69:0], callResR126);
  assign res = callResR126;
endmodule

module zdLLzilambda15200 (input logic [69:0] arg0,
  input logic [69:0] arg1,
  output logic [77:0] res);
  logic [69:0] gMainzir0;
  logic [69:0] gzdLLzicase16043;
  assign gMainzir0 = arg0;
  assign gzdLLzicase16043 = gMainzir0[69:0];
  assign res = {gzdLLzicase16043[69:62], arg1};
endmodule

module zdLLzilambda15411 (input logic [69:0] arg0,
  input logic [69:0] arg1,
  output logic [77:0] res);
  logic [69:0] gMainzir1;
  logic [69:0] gzdLLzicase16051;
  assign gMainzir1 = arg0;
  assign gzdLLzicase16051 = gMainzir1[69:0];
  assign res = {gzdLLzicase16051[61:54], arg1};
endmodule

module zdLLzilambda15413 (input logic [69:0] arg0,
  input logic [69:0] arg1,
  output logic [77:0] res);
  logic [69:0] gMainzir2;
  logic [69:0] gzdLLzicase16059;
  assign gMainzir2 = arg0;
  assign gzdLLzicase16059 = gMainzir2[69:0];
  assign res = {gzdLLzicase16059[53:46], arg1};
endmodule

module zdLLzilambda15415 (input logic [69:0] arg0,
  input logic [69:0] arg1,
  output logic [77:0] res);
  logic [69:0] gMainzir3;
  logic [69:0] gzdLLzicase16067;
  assign gMainzir3 = arg0;
  assign gzdLLzicase16067 = gMainzir3[69:0];
  assign res = {gzdLLzicase16067[45:38], arg1};
endmodule

module Mainziinputs (input logic [69:0] arg0,
  output logic [16:0] res);
  logic [69:0] gzdLLzicase14722;
  assign gzdLLzicase14722 = arg0;
  assign res = gzdLLzicase14722[31:15];
endmodule

module Mainzioutputs (input logic [69:0] arg0,
  output logic [14:0] res);
  logic [69:0] gzdLLzicase15902;
  assign gzdLLzicase15902 = arg0;
  assign res = gzdLLzicase15902[14:0];
endmodule

module Mainzipc (input logic [69:0] arg0,
  output logic [5:0] res);
  logic [69:0] gzdLLzicase15910;
  assign gzdLLzicase15910 = arg0;
  assign res = gzdLLzicase15910[37:32];
endmodule