module top_level (input logic [1:0] __in0,
  output logic [1:0] __out0);
  assign __out0 = 2'h1;
endmodule