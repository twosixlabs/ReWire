module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [63:0] __in0,
  input logic [63:0] __in1,
  output logic [63:0] __out0,
  output logic [63:0] __out1);
  logic [127:0] main_loop1_in;
  logic [127:0] main_compute1_in;
  logic [127:0] zll_main_compute_in;
  logic [130:0] zll_main_compute60_in;
  logic [7:0] zll_main_compute60_out;
  logic [130:0] zll_main_compute60_inR1;
  logic [7:0] zll_main_compute60_outR1;
  logic [130:0] zll_main_compute60_inR2;
  logic [7:0] zll_main_compute60_outR2;
  logic [130:0] zll_main_compute60_inR3;
  logic [7:0] zll_main_compute60_outR3;
  logic [130:0] zll_main_compute60_inR4;
  logic [7:0] zll_main_compute60_outR4;
  logic [130:0] zll_main_compute60_inR5;
  logic [7:0] zll_main_compute60_outR5;
  logic [130:0] zll_main_compute60_inR6;
  logic [7:0] zll_main_compute60_outR6;
  logic [130:0] zll_main_compute60_inR7;
  logic [7:0] zll_main_compute60_outR7;
  logic [130:0] zll_main_compute34_in;
  logic [7:0] zll_main_compute34_out;
  logic [130:0] zll_main_compute34_inR1;
  logic [7:0] zll_main_compute34_outR1;
  logic [130:0] zll_main_compute34_inR2;
  logic [7:0] zll_main_compute34_outR2;
  logic [130:0] zll_main_compute34_inR3;
  logic [7:0] zll_main_compute34_outR3;
  logic [130:0] zll_main_compute34_inR4;
  logic [7:0] zll_main_compute34_outR4;
  logic [130:0] zll_main_compute34_inR5;
  logic [7:0] zll_main_compute34_outR5;
  logic [130:0] zll_main_compute34_inR6;
  logic [7:0] zll_main_compute34_outR6;
  logic [130:0] zll_main_compute34_inR7;
  logic [7:0] zll_main_compute34_outR7;
  logic [128:0] zll_main_loop3_in;
  logic [128:0] zll_main_loop2_in;
  logic [0:0] __continue;
  logic [127:0] __resumption_tag;
  logic [127:0] __resumption_tag_next;
  assign main_loop1_in = __resumption_tag;
  assign main_compute1_in = main_loop1_in[127:0];
  assign zll_main_compute_in = main_compute1_in[127:0];
  assign zll_main_compute60_in = {zll_main_compute_in[127:64], zll_main_compute_in[63:0], 3'h0};
  ZLL_Main_compute60  inst (zll_main_compute60_in[130:67], zll_main_compute60_in[66:3], zll_main_compute60_in[2:0], zll_main_compute60_out);
  assign zll_main_compute60_inR1 = {zll_main_compute_in[127:64], zll_main_compute_in[63:0], 3'h1};
  ZLL_Main_compute60  instR1 (zll_main_compute60_inR1[130:67], zll_main_compute60_inR1[66:3], zll_main_compute60_inR1[2:0], zll_main_compute60_outR1);
  assign zll_main_compute60_inR2 = {zll_main_compute_in[127:64], zll_main_compute_in[63:0], 3'h2};
  ZLL_Main_compute60  instR2 (zll_main_compute60_inR2[130:67], zll_main_compute60_inR2[66:3], zll_main_compute60_inR2[2:0], zll_main_compute60_outR2);
  assign zll_main_compute60_inR3 = {zll_main_compute_in[127:64], zll_main_compute_in[63:0], 3'h3};
  ZLL_Main_compute60  instR3 (zll_main_compute60_inR3[130:67], zll_main_compute60_inR3[66:3], zll_main_compute60_inR3[2:0], zll_main_compute60_outR3);
  assign zll_main_compute60_inR4 = {zll_main_compute_in[127:64], zll_main_compute_in[63:0], 3'h4};
  ZLL_Main_compute60  instR4 (zll_main_compute60_inR4[130:67], zll_main_compute60_inR4[66:3], zll_main_compute60_inR4[2:0], zll_main_compute60_outR4);
  assign zll_main_compute60_inR5 = {zll_main_compute_in[127:64], zll_main_compute_in[63:0], 3'h5};
  ZLL_Main_compute60  instR5 (zll_main_compute60_inR5[130:67], zll_main_compute60_inR5[66:3], zll_main_compute60_inR5[2:0], zll_main_compute60_outR5);
  assign zll_main_compute60_inR6 = {zll_main_compute_in[127:64], zll_main_compute_in[63:0], 3'h6};
  ZLL_Main_compute60  instR6 (zll_main_compute60_inR6[130:67], zll_main_compute60_inR6[66:3], zll_main_compute60_inR6[2:0], zll_main_compute60_outR6);
  assign zll_main_compute60_inR7 = {zll_main_compute_in[127:64], zll_main_compute_in[63:0], 3'h7};
  ZLL_Main_compute60  instR7 (zll_main_compute60_inR7[130:67], zll_main_compute60_inR7[66:3], zll_main_compute60_inR7[2:0], zll_main_compute60_outR7);
  assign zll_main_compute34_in = {zll_main_compute_in[127:64], zll_main_compute_in[63:0], 3'h0};
  ZLL_Main_compute34  instR8 (zll_main_compute34_in[130:67], zll_main_compute34_in[66:3], zll_main_compute34_in[2:0], zll_main_compute34_out);
  assign zll_main_compute34_inR1 = {zll_main_compute_in[127:64], zll_main_compute_in[63:0], 3'h1};
  ZLL_Main_compute34  instR9 (zll_main_compute34_inR1[130:67], zll_main_compute34_inR1[66:3], zll_main_compute34_inR1[2:0], zll_main_compute34_outR1);
  assign zll_main_compute34_inR2 = {zll_main_compute_in[127:64], zll_main_compute_in[63:0], 3'h2};
  ZLL_Main_compute34  instR10 (zll_main_compute34_inR2[130:67], zll_main_compute34_inR2[66:3], zll_main_compute34_inR2[2:0], zll_main_compute34_outR2);
  assign zll_main_compute34_inR3 = {zll_main_compute_in[127:64], zll_main_compute_in[63:0], 3'h3};
  ZLL_Main_compute34  instR11 (zll_main_compute34_inR3[130:67], zll_main_compute34_inR3[66:3], zll_main_compute34_inR3[2:0], zll_main_compute34_outR3);
  assign zll_main_compute34_inR4 = {zll_main_compute_in[127:64], zll_main_compute_in[63:0], 3'h4};
  ZLL_Main_compute34  instR12 (zll_main_compute34_inR4[130:67], zll_main_compute34_inR4[66:3], zll_main_compute34_inR4[2:0], zll_main_compute34_outR4);
  assign zll_main_compute34_inR5 = {zll_main_compute_in[127:64], zll_main_compute_in[63:0], 3'h5};
  ZLL_Main_compute34  instR13 (zll_main_compute34_inR5[130:67], zll_main_compute34_inR5[66:3], zll_main_compute34_inR5[2:0], zll_main_compute34_outR5);
  assign zll_main_compute34_inR6 = {zll_main_compute_in[127:64], zll_main_compute_in[63:0], 3'h6};
  ZLL_Main_compute34  instR14 (zll_main_compute34_inR6[130:67], zll_main_compute34_inR6[66:3], zll_main_compute34_inR6[2:0], zll_main_compute34_outR6);
  assign zll_main_compute34_inR7 = {zll_main_compute_in[127:64], zll_main_compute_in[63:0], 3'h7};
  ZLL_Main_compute34  instR15 (zll_main_compute34_inR7[130:67], zll_main_compute34_inR7[66:3], zll_main_compute34_inR7[2:0], zll_main_compute34_outR7);
  assign zll_main_loop3_in = {1'h0, {zll_main_compute60_out, zll_main_compute60_outR1, zll_main_compute60_outR2, zll_main_compute60_outR3, zll_main_compute60_outR4, zll_main_compute60_outR5, zll_main_compute60_outR6, zll_main_compute60_outR7, zll_main_compute34_out, zll_main_compute34_outR1, zll_main_compute34_outR2, zll_main_compute34_outR3, zll_main_compute34_outR4, zll_main_compute34_outR5, zll_main_compute34_outR6, zll_main_compute34_outR7}};
  assign zll_main_loop2_in = zll_main_loop3_in[128:0];
  assign {__continue, __out0, __out1, __resumption_tag_next} = {1'h1, zll_main_loop2_in[127:0]};
  initial __resumption_tag <= {8'h80{1'h0}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      __resumption_tag <= {8'h80{1'h0}};
    end else begin
      __resumption_tag <= __resumption_tag_next;
    end
  end
endmodule

module ZLL_Main_compute72 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [255:0] binop_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [131:0] zll_main_compute66_in;
  logic [130:0] zll_main_compute43_in;
  logic [7:0] zll_main_compute43_out;
  logic [130:0] zll_main_compute43_inR1;
  logic [7:0] zll_main_compute43_outR1;
  logic [130:0] zll_main_compute43_inR2;
  logic [7:0] zll_main_compute43_outR2;
  logic [130:0] zll_main_compute43_inR3;
  logic [7:0] zll_main_compute43_outR3;
  logic [130:0] zll_main_compute43_inR4;
  logic [7:0] zll_main_compute43_outR4;
  logic [130:0] zll_main_compute43_inR5;
  logic [7:0] zll_main_compute43_outR5;
  logic [130:0] zll_main_compute43_inR6;
  logic [7:0] zll_main_compute43_outR6;
  logic [130:0] zll_main_compute43_inR7;
  logic [7:0] zll_main_compute43_outR7;
  logic [63:0] resize_inR2;
  logic [2:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR8;
  logic [2:0] resize_inR9;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR10;
  logic [131:0] zll_main_compute69_in;
  logic [130:0] zll_main_compute53_in;
  logic [7:0] zll_main_compute53_out;
  logic [130:0] zll_main_compute53_inR1;
  logic [7:0] zll_main_compute53_outR1;
  logic [130:0] zll_main_compute53_inR2;
  logic [7:0] zll_main_compute53_outR2;
  logic [130:0] zll_main_compute53_inR3;
  logic [7:0] zll_main_compute53_outR3;
  logic [130:0] zll_main_compute53_inR4;
  logic [7:0] zll_main_compute53_outR4;
  logic [130:0] zll_main_compute53_inR5;
  logic [7:0] zll_main_compute53_outR5;
  logic [130:0] zll_main_compute53_inR6;
  logic [7:0] zll_main_compute53_outR6;
  logic [130:0] zll_main_compute53_inR7;
  logic [7:0] zll_main_compute53_outR7;
  logic [63:0] resize_inR11;
  logic [2:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [127:0] resize_inR13;
  logic [2:0] resize_inR14;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR15;
  logic [2:0] resize_inR16;
  logic [255:0] binop_inR16;
  logic [255:0] binop_inR17;
  logic [255:0] binop_inR18;
  logic [255:0] binop_inR19;
  logic [127:0] resize_inR17;
  assign resize_in = arg2;
  assign binop_in = {128'(resize_in[2:0]), 128'h3};
  assign resize_inR1 = arg2;
  assign binop_inR1 = {128'(resize_inR1[2:0]), 128'h3};
  assign zll_main_compute66_in = {arg0, arg1, arg2, binop_inR1[255:128] < binop_inR1[127:0]};
  assign zll_main_compute43_in = {zll_main_compute66_in[131:68], zll_main_compute66_in[67:4], 3'h0};
  ZLL_Main_compute43  inst (zll_main_compute43_in[130:67], zll_main_compute43_in[66:3], zll_main_compute43_in[2:0], zll_main_compute43_out);
  assign zll_main_compute43_inR1 = {zll_main_compute66_in[131:68], zll_main_compute66_in[67:4], 3'h1};
  ZLL_Main_compute43  instR1 (zll_main_compute43_inR1[130:67], zll_main_compute43_inR1[66:3], zll_main_compute43_inR1[2:0], zll_main_compute43_outR1);
  assign zll_main_compute43_inR2 = {zll_main_compute66_in[131:68], zll_main_compute66_in[67:4], 3'h2};
  ZLL_Main_compute43  instR2 (zll_main_compute43_inR2[130:67], zll_main_compute43_inR2[66:3], zll_main_compute43_inR2[2:0], zll_main_compute43_outR2);
  assign zll_main_compute43_inR3 = {zll_main_compute66_in[131:68], zll_main_compute66_in[67:4], 3'h3};
  ZLL_Main_compute43  instR3 (zll_main_compute43_inR3[130:67], zll_main_compute43_inR3[66:3], zll_main_compute43_inR3[2:0], zll_main_compute43_outR3);
  assign zll_main_compute43_inR4 = {zll_main_compute66_in[131:68], zll_main_compute66_in[67:4], 3'h4};
  ZLL_Main_compute43  instR4 (zll_main_compute43_inR4[130:67], zll_main_compute43_inR4[66:3], zll_main_compute43_inR4[2:0], zll_main_compute43_outR4);
  assign zll_main_compute43_inR5 = {zll_main_compute66_in[131:68], zll_main_compute66_in[67:4], 3'h5};
  ZLL_Main_compute43  instR5 (zll_main_compute43_inR5[130:67], zll_main_compute43_inR5[66:3], zll_main_compute43_inR5[2:0], zll_main_compute43_outR5);
  assign zll_main_compute43_inR6 = {zll_main_compute66_in[131:68], zll_main_compute66_in[67:4], 3'h6};
  ZLL_Main_compute43  instR6 (zll_main_compute43_inR6[130:67], zll_main_compute43_inR6[66:3], zll_main_compute43_inR6[2:0], zll_main_compute43_outR6);
  assign zll_main_compute43_inR7 = {zll_main_compute66_in[131:68], zll_main_compute66_in[67:4], 3'h7};
  ZLL_Main_compute43  instR7 (zll_main_compute43_inR7[130:67], zll_main_compute43_inR7[66:3], zll_main_compute43_inR7[2:0], zll_main_compute43_outR7);
  assign resize_inR2 = {zll_main_compute43_out, zll_main_compute43_outR1, zll_main_compute43_outR2, zll_main_compute43_outR3, zll_main_compute43_outR4, zll_main_compute43_outR5, zll_main_compute43_outR6, zll_main_compute43_outR7};
  assign resize_inR3 = zll_main_compute66_in[3:1];
  assign binop_inR2 = {128'(resize_inR3[2:0]), 128'h3};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h8};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[2:0];
  assign binop_inR4 = {128'(resize_inR5[2:0]), 128'h2};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h8};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR6 = {128'(resize_inR7[2:0]), 128'h1};
  assign binop_inR7 = {binop_inR6[255:128] + binop_inR6[127:0], 128'h8};
  assign resize_inR8 = binop_inR7[255:128] % binop_inR7[127:0];
  assign resize_inR9 = resize_inR8[2:0];
  assign binop_inR8 = {128'h8, 128'(resize_inR9[2:0])};
  assign binop_inR9 = {binop_inR8[255:128] - binop_inR8[127:0], 128'h1};
  assign binop_inR10 = {binop_inR9[255:128] - binop_inR9[127:0], 128'h8};
  assign binop_inR11 = {128'(resize_inR2[63:0]), binop_inR10[255:128] * binop_inR10[127:0]};
  assign resize_inR10 = binop_inR11[255:128] >> binop_inR11[127:0];
  assign zll_main_compute69_in = {arg0, arg1, arg2, binop_in[255:128] < binop_in[127:0]};
  assign zll_main_compute53_in = {zll_main_compute69_in[131:68], zll_main_compute69_in[67:4], 3'h0};
  ZLL_Main_compute53  instR8 (zll_main_compute53_in[130:67], zll_main_compute53_in[66:3], zll_main_compute53_in[2:0], zll_main_compute53_out);
  assign zll_main_compute53_inR1 = {zll_main_compute69_in[131:68], zll_main_compute69_in[67:4], 3'h1};
  ZLL_Main_compute53  instR9 (zll_main_compute53_inR1[130:67], zll_main_compute53_inR1[66:3], zll_main_compute53_inR1[2:0], zll_main_compute53_outR1);
  assign zll_main_compute53_inR2 = {zll_main_compute69_in[131:68], zll_main_compute69_in[67:4], 3'h2};
  ZLL_Main_compute53  instR10 (zll_main_compute53_inR2[130:67], zll_main_compute53_inR2[66:3], zll_main_compute53_inR2[2:0], zll_main_compute53_outR2);
  assign zll_main_compute53_inR3 = {zll_main_compute69_in[131:68], zll_main_compute69_in[67:4], 3'h3};
  ZLL_Main_compute53  instR11 (zll_main_compute53_inR3[130:67], zll_main_compute53_inR3[66:3], zll_main_compute53_inR3[2:0], zll_main_compute53_outR3);
  assign zll_main_compute53_inR4 = {zll_main_compute69_in[131:68], zll_main_compute69_in[67:4], 3'h4};
  ZLL_Main_compute53  instR12 (zll_main_compute53_inR4[130:67], zll_main_compute53_inR4[66:3], zll_main_compute53_inR4[2:0], zll_main_compute53_outR4);
  assign zll_main_compute53_inR5 = {zll_main_compute69_in[131:68], zll_main_compute69_in[67:4], 3'h5};
  ZLL_Main_compute53  instR13 (zll_main_compute53_inR5[130:67], zll_main_compute53_inR5[66:3], zll_main_compute53_inR5[2:0], zll_main_compute53_outR5);
  assign zll_main_compute53_inR6 = {zll_main_compute69_in[131:68], zll_main_compute69_in[67:4], 3'h6};
  ZLL_Main_compute53  instR14 (zll_main_compute53_inR6[130:67], zll_main_compute53_inR6[66:3], zll_main_compute53_inR6[2:0], zll_main_compute53_outR6);
  assign zll_main_compute53_inR7 = {zll_main_compute69_in[131:68], zll_main_compute69_in[67:4], 3'h7};
  ZLL_Main_compute53  instR15 (zll_main_compute53_inR7[130:67], zll_main_compute53_inR7[66:3], zll_main_compute53_inR7[2:0], zll_main_compute53_outR7);
  assign resize_inR11 = {zll_main_compute53_out, zll_main_compute53_outR1, zll_main_compute53_outR2, zll_main_compute53_outR3, zll_main_compute53_outR4, zll_main_compute53_outR5, zll_main_compute53_outR6, zll_main_compute53_outR7};
  assign resize_inR12 = zll_main_compute69_in[3:1];
  assign binop_inR12 = {128'(resize_inR12[2:0]), 128'h2};
  assign binop_inR13 = {binop_inR12[255:128] * binop_inR12[127:0], 128'h8};
  assign resize_inR13 = binop_inR13[255:128] % binop_inR13[127:0];
  assign resize_inR14 = resize_inR13[2:0];
  assign binop_inR14 = {128'(resize_inR14[2:0]), 128'h1};
  assign binop_inR15 = {binop_inR14[255:128] + binop_inR14[127:0], 128'h8};
  assign resize_inR15 = binop_inR15[255:128] % binop_inR15[127:0];
  assign resize_inR16 = resize_inR15[2:0];
  assign binop_inR16 = {128'h8, 128'(resize_inR16[2:0])};
  assign binop_inR17 = {binop_inR16[255:128] - binop_inR16[127:0], 128'h1};
  assign binop_inR18 = {binop_inR17[255:128] - binop_inR17[127:0], 128'h8};
  assign binop_inR19 = {128'(resize_inR11[63:0]), binop_inR18[255:128] * binop_inR18[127:0]};
  assign resize_inR17 = binop_inR19[255:128] >> binop_inR19[127:0];
  assign res = (zll_main_compute69_in[0] == 1'h1) ? resize_inR17[7:0] : resize_inR10[7:0];
endmodule

module ZLL_Main_compute65 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [255:0] binop_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [131:0] zll_main_compute41_in;
  logic [130:0] zll_main_compute37_in;
  logic [7:0] zll_main_compute37_out;
  logic [130:0] zll_main_compute37_inR1;
  logic [7:0] zll_main_compute37_outR1;
  logic [130:0] zll_main_compute37_inR2;
  logic [7:0] zll_main_compute37_outR2;
  logic [130:0] zll_main_compute37_inR3;
  logic [7:0] zll_main_compute37_outR3;
  logic [130:0] zll_main_compute37_inR4;
  logic [7:0] zll_main_compute37_outR4;
  logic [130:0] zll_main_compute37_inR5;
  logic [7:0] zll_main_compute37_outR5;
  logic [130:0] zll_main_compute37_inR6;
  logic [7:0] zll_main_compute37_outR6;
  logic [130:0] zll_main_compute37_inR7;
  logic [7:0] zll_main_compute37_outR7;
  logic [63:0] resize_inR2;
  logic [2:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR8;
  logic [131:0] zll_main_compute42_in;
  logic [130:0] zll_main_compute53_in;
  logic [7:0] zll_main_compute53_out;
  logic [130:0] zll_main_compute53_inR1;
  logic [7:0] zll_main_compute53_outR1;
  logic [130:0] zll_main_compute53_inR2;
  logic [7:0] zll_main_compute53_outR2;
  logic [130:0] zll_main_compute53_inR3;
  logic [7:0] zll_main_compute53_outR3;
  logic [130:0] zll_main_compute53_inR4;
  logic [7:0] zll_main_compute53_outR4;
  logic [130:0] zll_main_compute53_inR5;
  logic [7:0] zll_main_compute53_outR5;
  logic [130:0] zll_main_compute53_inR6;
  logic [7:0] zll_main_compute53_outR6;
  logic [130:0] zll_main_compute53_inR7;
  logic [7:0] zll_main_compute53_outR7;
  logic [63:0] resize_inR9;
  logic [2:0] resize_inR10;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR11;
  logic [2:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR13;
  assign resize_in = arg2;
  assign binop_in = {128'(resize_in[2:0]), 128'h3};
  assign resize_inR1 = arg2;
  assign binop_inR1 = {128'(resize_inR1[2:0]), 128'h3};
  assign zll_main_compute41_in = {arg0, arg1, arg2, binop_inR1[255:128] < binop_inR1[127:0]};
  assign zll_main_compute37_in = {zll_main_compute41_in[131:68], zll_main_compute41_in[67:4], 3'h0};
  ZLL_Main_compute37  inst (zll_main_compute37_in[130:67], zll_main_compute37_in[66:3], zll_main_compute37_in[2:0], zll_main_compute37_out);
  assign zll_main_compute37_inR1 = {zll_main_compute41_in[131:68], zll_main_compute41_in[67:4], 3'h1};
  ZLL_Main_compute37  instR1 (zll_main_compute37_inR1[130:67], zll_main_compute37_inR1[66:3], zll_main_compute37_inR1[2:0], zll_main_compute37_outR1);
  assign zll_main_compute37_inR2 = {zll_main_compute41_in[131:68], zll_main_compute41_in[67:4], 3'h2};
  ZLL_Main_compute37  instR2 (zll_main_compute37_inR2[130:67], zll_main_compute37_inR2[66:3], zll_main_compute37_inR2[2:0], zll_main_compute37_outR2);
  assign zll_main_compute37_inR3 = {zll_main_compute41_in[131:68], zll_main_compute41_in[67:4], 3'h3};
  ZLL_Main_compute37  instR3 (zll_main_compute37_inR3[130:67], zll_main_compute37_inR3[66:3], zll_main_compute37_inR3[2:0], zll_main_compute37_outR3);
  assign zll_main_compute37_inR4 = {zll_main_compute41_in[131:68], zll_main_compute41_in[67:4], 3'h4};
  ZLL_Main_compute37  instR4 (zll_main_compute37_inR4[130:67], zll_main_compute37_inR4[66:3], zll_main_compute37_inR4[2:0], zll_main_compute37_outR4);
  assign zll_main_compute37_inR5 = {zll_main_compute41_in[131:68], zll_main_compute41_in[67:4], 3'h5};
  ZLL_Main_compute37  instR5 (zll_main_compute37_inR5[130:67], zll_main_compute37_inR5[66:3], zll_main_compute37_inR5[2:0], zll_main_compute37_outR5);
  assign zll_main_compute37_inR6 = {zll_main_compute41_in[131:68], zll_main_compute41_in[67:4], 3'h6};
  ZLL_Main_compute37  instR6 (zll_main_compute37_inR6[130:67], zll_main_compute37_inR6[66:3], zll_main_compute37_inR6[2:0], zll_main_compute37_outR6);
  assign zll_main_compute37_inR7 = {zll_main_compute41_in[131:68], zll_main_compute41_in[67:4], 3'h7};
  ZLL_Main_compute37  instR7 (zll_main_compute37_inR7[130:67], zll_main_compute37_inR7[66:3], zll_main_compute37_inR7[2:0], zll_main_compute37_outR7);
  assign resize_inR2 = {zll_main_compute37_out, zll_main_compute37_outR1, zll_main_compute37_outR2, zll_main_compute37_outR3, zll_main_compute37_outR4, zll_main_compute37_outR5, zll_main_compute37_outR6, zll_main_compute37_outR7};
  assign resize_inR3 = zll_main_compute41_in[3:1];
  assign binop_inR2 = {128'(resize_inR3[2:0]), 128'h3};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h8};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[2:0];
  assign binop_inR4 = {128'(resize_inR5[2:0]), 128'h2};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h8};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR6 = {128'h8, 128'(resize_inR7[2:0])};
  assign binop_inR7 = {binop_inR6[255:128] - binop_inR6[127:0], 128'h1};
  assign binop_inR8 = {binop_inR7[255:128] - binop_inR7[127:0], 128'h8};
  assign binop_inR9 = {128'(resize_inR2[63:0]), binop_inR8[255:128] * binop_inR8[127:0]};
  assign resize_inR8 = binop_inR9[255:128] >> binop_inR9[127:0];
  assign zll_main_compute42_in = {arg0, arg1, arg2, binop_in[255:128] < binop_in[127:0]};
  assign zll_main_compute53_in = {zll_main_compute42_in[131:68], zll_main_compute42_in[67:4], 3'h0};
  ZLL_Main_compute53  instR8 (zll_main_compute53_in[130:67], zll_main_compute53_in[66:3], zll_main_compute53_in[2:0], zll_main_compute53_out);
  assign zll_main_compute53_inR1 = {zll_main_compute42_in[131:68], zll_main_compute42_in[67:4], 3'h1};
  ZLL_Main_compute53  instR9 (zll_main_compute53_inR1[130:67], zll_main_compute53_inR1[66:3], zll_main_compute53_inR1[2:0], zll_main_compute53_outR1);
  assign zll_main_compute53_inR2 = {zll_main_compute42_in[131:68], zll_main_compute42_in[67:4], 3'h2};
  ZLL_Main_compute53  instR10 (zll_main_compute53_inR2[130:67], zll_main_compute53_inR2[66:3], zll_main_compute53_inR2[2:0], zll_main_compute53_outR2);
  assign zll_main_compute53_inR3 = {zll_main_compute42_in[131:68], zll_main_compute42_in[67:4], 3'h3};
  ZLL_Main_compute53  instR11 (zll_main_compute53_inR3[130:67], zll_main_compute53_inR3[66:3], zll_main_compute53_inR3[2:0], zll_main_compute53_outR3);
  assign zll_main_compute53_inR4 = {zll_main_compute42_in[131:68], zll_main_compute42_in[67:4], 3'h4};
  ZLL_Main_compute53  instR12 (zll_main_compute53_inR4[130:67], zll_main_compute53_inR4[66:3], zll_main_compute53_inR4[2:0], zll_main_compute53_outR4);
  assign zll_main_compute53_inR5 = {zll_main_compute42_in[131:68], zll_main_compute42_in[67:4], 3'h5};
  ZLL_Main_compute53  instR13 (zll_main_compute53_inR5[130:67], zll_main_compute53_inR5[66:3], zll_main_compute53_inR5[2:0], zll_main_compute53_outR5);
  assign zll_main_compute53_inR6 = {zll_main_compute42_in[131:68], zll_main_compute42_in[67:4], 3'h6};
  ZLL_Main_compute53  instR14 (zll_main_compute53_inR6[130:67], zll_main_compute53_inR6[66:3], zll_main_compute53_inR6[2:0], zll_main_compute53_outR6);
  assign zll_main_compute53_inR7 = {zll_main_compute42_in[131:68], zll_main_compute42_in[67:4], 3'h7};
  ZLL_Main_compute53  instR15 (zll_main_compute53_inR7[130:67], zll_main_compute53_inR7[66:3], zll_main_compute53_inR7[2:0], zll_main_compute53_outR7);
  assign resize_inR9 = {zll_main_compute53_out, zll_main_compute53_outR1, zll_main_compute53_outR2, zll_main_compute53_outR3, zll_main_compute53_outR4, zll_main_compute53_outR5, zll_main_compute53_outR6, zll_main_compute53_outR7};
  assign resize_inR10 = zll_main_compute42_in[3:1];
  assign binop_inR10 = {128'(resize_inR10[2:0]), 128'h2};
  assign binop_inR11 = {binop_inR10[255:128] * binop_inR10[127:0], 128'h8};
  assign resize_inR11 = binop_inR11[255:128] % binop_inR11[127:0];
  assign resize_inR12 = resize_inR11[2:0];
  assign binop_inR12 = {128'h8, 128'(resize_inR12[2:0])};
  assign binop_inR13 = {binop_inR12[255:128] - binop_inR12[127:0], 128'h1};
  assign binop_inR14 = {binop_inR13[255:128] - binop_inR13[127:0], 128'h8};
  assign binop_inR15 = {128'(resize_inR9[63:0]), binop_inR14[255:128] * binop_inR14[127:0]};
  assign resize_inR13 = binop_inR15[255:128] >> binop_inR15[127:0];
  assign res = (zll_main_compute42_in[0] == 1'h1) ? resize_inR13[7:0] : resize_inR8[7:0];
endmodule

module ReWire_Prelude_not (input logic [0:0] arg0,
  output logic [0:0] res);
  logic [0:0] lit_in;
  assign lit_in = arg0;
  assign res = (lit_in[0] == 1'h1) ? 1'h0 : 1'h1;
endmodule

module ZLL_Main_compute60 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [127:0] resize_inR1;
  logic [0:0] msbit_in;
  logic [0:0] rewire_prelude_not_in;
  logic [0:0] rewire_prelude_not_out;
  logic [2:0] resize_inR2;
  logic [127:0] resize_inR3;
  logic [0:0] msbit_inR1;
  logic [0:0] rewire_prelude_not_inR1;
  logic [0:0] rewire_prelude_not_outR1;
  logic [131:0] zll_main_compute26_in;
  logic [130:0] zll_main_compute72_in;
  logic [7:0] zll_main_compute72_out;
  logic [130:0] zll_main_compute72_inR1;
  logic [7:0] zll_main_compute72_outR1;
  logic [130:0] zll_main_compute72_inR2;
  logic [7:0] zll_main_compute72_outR2;
  logic [130:0] zll_main_compute72_inR3;
  logic [7:0] zll_main_compute72_outR3;
  logic [130:0] zll_main_compute72_inR4;
  logic [7:0] zll_main_compute72_outR4;
  logic [130:0] zll_main_compute72_inR5;
  logic [7:0] zll_main_compute72_outR5;
  logic [130:0] zll_main_compute72_inR6;
  logic [7:0] zll_main_compute72_outR6;
  logic [130:0] zll_main_compute72_inR7;
  logic [7:0] zll_main_compute72_outR7;
  logic [63:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR8;
  logic [2:0] resize_inR9;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR10;
  logic [131:0] zll_main_compute15_in;
  logic [130:0] zll_main_compute65_in;
  logic [7:0] zll_main_compute65_out;
  logic [130:0] zll_main_compute65_inR1;
  logic [7:0] zll_main_compute65_outR1;
  logic [130:0] zll_main_compute65_inR2;
  logic [7:0] zll_main_compute65_outR2;
  logic [130:0] zll_main_compute65_inR3;
  logic [7:0] zll_main_compute65_outR3;
  logic [130:0] zll_main_compute65_inR4;
  logic [7:0] zll_main_compute65_outR4;
  logic [130:0] zll_main_compute65_inR5;
  logic [7:0] zll_main_compute65_outR5;
  logic [130:0] zll_main_compute65_inR6;
  logic [7:0] zll_main_compute65_outR6;
  logic [130:0] zll_main_compute65_inR7;
  logic [7:0] zll_main_compute65_outR7;
  logic [63:0] resize_inR11;
  logic [2:0] resize_inR12;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR13;
  logic [2:0] resize_inR14;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [127:0] resize_inR15;
  assign resize_in = arg2;
  assign resize_inR1 = 128'(resize_in[2:0]);
  assign msbit_in = resize_inR1[0];
  assign rewire_prelude_not_in = msbit_in[0];
  ReWire_Prelude_not  inst (rewire_prelude_not_in[0], rewire_prelude_not_out);
  assign resize_inR2 = arg2;
  assign resize_inR3 = 128'(resize_inR2[2:0]);
  assign msbit_inR1 = resize_inR3[0];
  assign rewire_prelude_not_inR1 = msbit_inR1[0];
  ReWire_Prelude_not  instR1 (rewire_prelude_not_inR1[0], rewire_prelude_not_outR1);
  assign zll_main_compute26_in = {arg0, arg1, arg2, rewire_prelude_not_outR1};
  assign zll_main_compute72_in = {zll_main_compute26_in[131:68], zll_main_compute26_in[67:4], 3'h0};
  ZLL_Main_compute72  instR2 (zll_main_compute72_in[130:67], zll_main_compute72_in[66:3], zll_main_compute72_in[2:0], zll_main_compute72_out);
  assign zll_main_compute72_inR1 = {zll_main_compute26_in[131:68], zll_main_compute26_in[67:4], 3'h1};
  ZLL_Main_compute72  instR3 (zll_main_compute72_inR1[130:67], zll_main_compute72_inR1[66:3], zll_main_compute72_inR1[2:0], zll_main_compute72_outR1);
  assign zll_main_compute72_inR2 = {zll_main_compute26_in[131:68], zll_main_compute26_in[67:4], 3'h2};
  ZLL_Main_compute72  instR4 (zll_main_compute72_inR2[130:67], zll_main_compute72_inR2[66:3], zll_main_compute72_inR2[2:0], zll_main_compute72_outR2);
  assign zll_main_compute72_inR3 = {zll_main_compute26_in[131:68], zll_main_compute26_in[67:4], 3'h3};
  ZLL_Main_compute72  instR5 (zll_main_compute72_inR3[130:67], zll_main_compute72_inR3[66:3], zll_main_compute72_inR3[2:0], zll_main_compute72_outR3);
  assign zll_main_compute72_inR4 = {zll_main_compute26_in[131:68], zll_main_compute26_in[67:4], 3'h4};
  ZLL_Main_compute72  instR6 (zll_main_compute72_inR4[130:67], zll_main_compute72_inR4[66:3], zll_main_compute72_inR4[2:0], zll_main_compute72_outR4);
  assign zll_main_compute72_inR5 = {zll_main_compute26_in[131:68], zll_main_compute26_in[67:4], 3'h5};
  ZLL_Main_compute72  instR7 (zll_main_compute72_inR5[130:67], zll_main_compute72_inR5[66:3], zll_main_compute72_inR5[2:0], zll_main_compute72_outR5);
  assign zll_main_compute72_inR6 = {zll_main_compute26_in[131:68], zll_main_compute26_in[67:4], 3'h6};
  ZLL_Main_compute72  instR8 (zll_main_compute72_inR6[130:67], zll_main_compute72_inR6[66:3], zll_main_compute72_inR6[2:0], zll_main_compute72_outR6);
  assign zll_main_compute72_inR7 = {zll_main_compute26_in[131:68], zll_main_compute26_in[67:4], 3'h7};
  ZLL_Main_compute72  instR9 (zll_main_compute72_inR7[130:67], zll_main_compute72_inR7[66:3], zll_main_compute72_inR7[2:0], zll_main_compute72_outR7);
  assign resize_inR4 = {zll_main_compute72_out, zll_main_compute72_outR1, zll_main_compute72_outR2, zll_main_compute72_outR3, zll_main_compute72_outR4, zll_main_compute72_outR5, zll_main_compute72_outR6, zll_main_compute72_outR7};
  assign resize_inR5 = zll_main_compute26_in[3:1];
  assign binop_in = {128'(resize_inR5[2:0]), 128'h1};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h8};
  assign resize_inR6 = binop_inR1[255:128] % binop_inR1[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR2 = {128'(resize_inR7[2:0]), 128'h2};
  assign binop_inR3 = {binop_inR2[255:128] / binop_inR2[127:0], 128'h8};
  assign resize_inR8 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR9 = resize_inR8[2:0];
  assign binop_inR4 = {128'h8, 128'(resize_inR9[2:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h8};
  assign binop_inR7 = {128'(resize_inR4[63:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR10 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign zll_main_compute15_in = {arg0, arg1, arg2, rewire_prelude_not_out};
  assign zll_main_compute65_in = {zll_main_compute15_in[131:68], zll_main_compute15_in[67:4], 3'h0};
  ZLL_Main_compute65  instR10 (zll_main_compute65_in[130:67], zll_main_compute65_in[66:3], zll_main_compute65_in[2:0], zll_main_compute65_out);
  assign zll_main_compute65_inR1 = {zll_main_compute15_in[131:68], zll_main_compute15_in[67:4], 3'h1};
  ZLL_Main_compute65  instR11 (zll_main_compute65_inR1[130:67], zll_main_compute65_inR1[66:3], zll_main_compute65_inR1[2:0], zll_main_compute65_outR1);
  assign zll_main_compute65_inR2 = {zll_main_compute15_in[131:68], zll_main_compute15_in[67:4], 3'h2};
  ZLL_Main_compute65  instR12 (zll_main_compute65_inR2[130:67], zll_main_compute65_inR2[66:3], zll_main_compute65_inR2[2:0], zll_main_compute65_outR2);
  assign zll_main_compute65_inR3 = {zll_main_compute15_in[131:68], zll_main_compute15_in[67:4], 3'h3};
  ZLL_Main_compute65  instR13 (zll_main_compute65_inR3[130:67], zll_main_compute65_inR3[66:3], zll_main_compute65_inR3[2:0], zll_main_compute65_outR3);
  assign zll_main_compute65_inR4 = {zll_main_compute15_in[131:68], zll_main_compute15_in[67:4], 3'h4};
  ZLL_Main_compute65  instR14 (zll_main_compute65_inR4[130:67], zll_main_compute65_inR4[66:3], zll_main_compute65_inR4[2:0], zll_main_compute65_outR4);
  assign zll_main_compute65_inR5 = {zll_main_compute15_in[131:68], zll_main_compute15_in[67:4], 3'h5};
  ZLL_Main_compute65  instR15 (zll_main_compute65_inR5[130:67], zll_main_compute65_inR5[66:3], zll_main_compute65_inR5[2:0], zll_main_compute65_outR5);
  assign zll_main_compute65_inR6 = {zll_main_compute15_in[131:68], zll_main_compute15_in[67:4], 3'h6};
  ZLL_Main_compute65  instR16 (zll_main_compute65_inR6[130:67], zll_main_compute65_inR6[66:3], zll_main_compute65_inR6[2:0], zll_main_compute65_outR6);
  assign zll_main_compute65_inR7 = {zll_main_compute15_in[131:68], zll_main_compute15_in[67:4], 3'h7};
  ZLL_Main_compute65  instR17 (zll_main_compute65_inR7[130:67], zll_main_compute65_inR7[66:3], zll_main_compute65_inR7[2:0], zll_main_compute65_outR7);
  assign resize_inR11 = {zll_main_compute65_out, zll_main_compute65_outR1, zll_main_compute65_outR2, zll_main_compute65_outR3, zll_main_compute65_outR4, zll_main_compute65_outR5, zll_main_compute65_outR6, zll_main_compute65_outR7};
  assign resize_inR12 = zll_main_compute15_in[3:1];
  assign binop_inR8 = {128'(resize_inR12[2:0]), 128'h2};
  assign binop_inR9 = {binop_inR8[255:128] / binop_inR8[127:0], 128'h8};
  assign resize_inR13 = binop_inR9[255:128] % binop_inR9[127:0];
  assign resize_inR14 = resize_inR13[2:0];
  assign binop_inR10 = {128'h8, 128'(resize_inR14[2:0])};
  assign binop_inR11 = {binop_inR10[255:128] - binop_inR10[127:0], 128'h1};
  assign binop_inR12 = {binop_inR11[255:128] - binop_inR11[127:0], 128'h8};
  assign binop_inR13 = {128'(resize_inR11[63:0]), binop_inR12[255:128] * binop_inR12[127:0]};
  assign resize_inR15 = binop_inR13[255:128] >> binop_inR13[127:0];
  assign res = (zll_main_compute15_in[0] == 1'h1) ? resize_inR15[7:0] : resize_inR10[7:0];
endmodule

module ZLL_Main_compute53 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [255:0] binop_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [67:0] zll_main_compute51_in;
  logic [63:0] resize_inR2;
  logic [2:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR8;
  logic [2:0] resize_inR9;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR10;
  logic [67:0] zll_main_compute71_in;
  logic [63:0] resize_inR11;
  logic [2:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [127:0] resize_inR13;
  logic [2:0] resize_inR14;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR15;
  logic [2:0] resize_inR16;
  logic [255:0] binop_inR16;
  logic [255:0] binop_inR17;
  logic [255:0] binop_inR18;
  logic [255:0] binop_inR19;
  logic [127:0] resize_inR17;
  assign resize_in = arg2;
  assign binop_in = {128'(resize_in[2:0]), 128'h3};
  assign resize_inR1 = arg2;
  assign binop_inR1 = {128'(resize_inR1[2:0]), 128'h3};
  assign zll_main_compute51_in = {arg1, arg2, binop_inR1[255:128] < binop_inR1[127:0]};
  assign resize_inR2 = zll_main_compute51_in[67:4];
  assign resize_inR3 = zll_main_compute51_in[3:1];
  assign binop_inR2 = {128'(resize_inR3[2:0]), 128'h3};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h8};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[2:0];
  assign binop_inR4 = {128'(resize_inR5[2:0]), 128'h2};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h8};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR6 = {128'(resize_inR7[2:0]), 128'h1};
  assign binop_inR7 = {binop_inR6[255:128] + binop_inR6[127:0], 128'h8};
  assign resize_inR8 = binop_inR7[255:128] % binop_inR7[127:0];
  assign resize_inR9 = resize_inR8[2:0];
  assign binop_inR8 = {128'h8, 128'(resize_inR9[2:0])};
  assign binop_inR9 = {binop_inR8[255:128] - binop_inR8[127:0], 128'h1};
  assign binop_inR10 = {binop_inR9[255:128] - binop_inR9[127:0], 128'h8};
  assign binop_inR11 = {128'(resize_inR2[63:0]), binop_inR10[255:128] * binop_inR10[127:0]};
  assign resize_inR10 = binop_inR11[255:128] >> binop_inR11[127:0];
  assign zll_main_compute71_in = {arg0, arg2, binop_in[255:128] < binop_in[127:0]};
  assign resize_inR11 = zll_main_compute71_in[67:4];
  assign resize_inR12 = zll_main_compute71_in[3:1];
  assign binop_inR12 = {128'(resize_inR12[2:0]), 128'h2};
  assign binop_inR13 = {binop_inR12[255:128] * binop_inR12[127:0], 128'h8};
  assign resize_inR13 = binop_inR13[255:128] % binop_inR13[127:0];
  assign resize_inR14 = resize_inR13[2:0];
  assign binop_inR14 = {128'(resize_inR14[2:0]), 128'h1};
  assign binop_inR15 = {binop_inR14[255:128] + binop_inR14[127:0], 128'h8};
  assign resize_inR15 = binop_inR15[255:128] % binop_inR15[127:0];
  assign resize_inR16 = resize_inR15[2:0];
  assign binop_inR16 = {128'h8, 128'(resize_inR16[2:0])};
  assign binop_inR17 = {binop_inR16[255:128] - binop_inR16[127:0], 128'h1};
  assign binop_inR18 = {binop_inR17[255:128] - binop_inR17[127:0], 128'h8};
  assign binop_inR19 = {128'(resize_inR11[63:0]), binop_inR18[255:128] * binop_inR18[127:0]};
  assign resize_inR17 = binop_inR19[255:128] >> binop_inR19[127:0];
  assign res = (zll_main_compute71_in[0] == 1'h1) ? resize_inR17[7:0] : resize_inR10[7:0];
endmodule

module ZLL_Main_compute43 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [255:0] binop_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [67:0] zll_main_compute48_in;
  logic [63:0] resize_inR2;
  logic [2:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR8;
  logic [67:0] zll_main_compute75_in;
  logic [63:0] resize_inR9;
  logic [2:0] resize_inR10;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR11;
  logic [2:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR13;
  assign resize_in = arg2;
  assign binop_in = {128'(resize_in[2:0]), 128'h3};
  assign resize_inR1 = arg2;
  assign binop_inR1 = {128'(resize_inR1[2:0]), 128'h3};
  assign zll_main_compute48_in = {arg1, arg2, binop_inR1[255:128] < binop_inR1[127:0]};
  assign resize_inR2 = zll_main_compute48_in[67:4];
  assign resize_inR3 = zll_main_compute48_in[3:1];
  assign binop_inR2 = {128'(resize_inR3[2:0]), 128'h3};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h8};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[2:0];
  assign binop_inR4 = {128'(resize_inR5[2:0]), 128'h2};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h8};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR6 = {128'h8, 128'(resize_inR7[2:0])};
  assign binop_inR7 = {binop_inR6[255:128] - binop_inR6[127:0], 128'h1};
  assign binop_inR8 = {binop_inR7[255:128] - binop_inR7[127:0], 128'h8};
  assign binop_inR9 = {128'(resize_inR2[63:0]), binop_inR8[255:128] * binop_inR8[127:0]};
  assign resize_inR8 = binop_inR9[255:128] >> binop_inR9[127:0];
  assign zll_main_compute75_in = {arg0, arg2, binop_in[255:128] < binop_in[127:0]};
  assign resize_inR9 = zll_main_compute75_in[67:4];
  assign resize_inR10 = zll_main_compute75_in[3:1];
  assign binop_inR10 = {128'(resize_inR10[2:0]), 128'h2};
  assign binop_inR11 = {binop_inR10[255:128] * binop_inR10[127:0], 128'h8};
  assign resize_inR11 = binop_inR11[255:128] % binop_inR11[127:0];
  assign resize_inR12 = resize_inR11[2:0];
  assign binop_inR12 = {128'h8, 128'(resize_inR12[2:0])};
  assign binop_inR13 = {binop_inR12[255:128] - binop_inR12[127:0], 128'h1};
  assign binop_inR14 = {binop_inR13[255:128] - binop_inR13[127:0], 128'h8};
  assign binop_inR15 = {128'(resize_inR9[63:0]), binop_inR14[255:128] * binop_inR14[127:0]};
  assign resize_inR13 = binop_inR15[255:128] >> binop_inR15[127:0];
  assign res = (zll_main_compute75_in[0] == 1'h1) ? resize_inR13[7:0] : resize_inR8[7:0];
endmodule

module ZLL_Main_compute37 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [255:0] binop_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [67:0] zll_main_compute78_in;
  logic [63:0] resize_inR2;
  logic [2:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR8;
  logic [67:0] zll_main_compute58_in;
  logic [63:0] resize_inR9;
  logic [2:0] resize_inR10;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR11;
  logic [2:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR13;
  assign resize_in = arg2;
  assign binop_in = {128'(resize_in[2:0]), 128'h3};
  assign resize_inR1 = arg2;
  assign binop_inR1 = {128'(resize_inR1[2:0]), 128'h3};
  assign zll_main_compute78_in = {arg2, arg1, binop_inR1[255:128] < binop_inR1[127:0]};
  assign resize_inR2 = zll_main_compute78_in[64:1];
  assign resize_inR3 = zll_main_compute78_in[67:65];
  assign binop_inR2 = {128'(resize_inR3[2:0]), 128'h3};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h8};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[2:0];
  assign binop_inR4 = {128'(resize_inR5[2:0]), 128'h2};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h8};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR6 = {128'h8, 128'(resize_inR7[2:0])};
  assign binop_inR7 = {binop_inR6[255:128] - binop_inR6[127:0], 128'h1};
  assign binop_inR8 = {binop_inR7[255:128] - binop_inR7[127:0], 128'h8};
  assign binop_inR9 = {128'(resize_inR2[63:0]), binop_inR8[255:128] * binop_inR8[127:0]};
  assign resize_inR8 = binop_inR9[255:128] >> binop_inR9[127:0];
  assign zll_main_compute58_in = {arg2, arg0, binop_in[255:128] < binop_in[127:0]};
  assign resize_inR9 = zll_main_compute58_in[64:1];
  assign resize_inR10 = zll_main_compute58_in[67:65];
  assign binop_inR10 = {128'(resize_inR10[2:0]), 128'h2};
  assign binop_inR11 = {binop_inR10[255:128] * binop_inR10[127:0], 128'h8};
  assign resize_inR11 = binop_inR11[255:128] % binop_inR11[127:0];
  assign resize_inR12 = resize_inR11[2:0];
  assign binop_inR12 = {128'h8, 128'(resize_inR12[2:0])};
  assign binop_inR13 = {binop_inR12[255:128] - binop_inR12[127:0], 128'h1};
  assign binop_inR14 = {binop_inR13[255:128] - binop_inR13[127:0], 128'h8};
  assign binop_inR15 = {128'(resize_inR9[63:0]), binop_inR14[255:128] * binop_inR14[127:0]};
  assign resize_inR13 = binop_inR15[255:128] >> binop_inR15[127:0];
  assign res = (zll_main_compute58_in[0] == 1'h1) ? resize_inR13[7:0] : resize_inR8[7:0];
endmodule

module ZLL_Main_compute36 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [255:0] binop_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [131:0] zll_main_compute59_in;
  logic [130:0] zll_main_compute43_in;
  logic [7:0] zll_main_compute43_out;
  logic [130:0] zll_main_compute43_inR1;
  logic [7:0] zll_main_compute43_outR1;
  logic [130:0] zll_main_compute43_inR2;
  logic [7:0] zll_main_compute43_outR2;
  logic [130:0] zll_main_compute43_inR3;
  logic [7:0] zll_main_compute43_outR3;
  logic [130:0] zll_main_compute43_inR4;
  logic [7:0] zll_main_compute43_outR4;
  logic [130:0] zll_main_compute43_inR5;
  logic [7:0] zll_main_compute43_outR5;
  logic [130:0] zll_main_compute43_inR6;
  logic [7:0] zll_main_compute43_outR6;
  logic [130:0] zll_main_compute43_inR7;
  logic [7:0] zll_main_compute43_outR7;
  logic [63:0] resize_inR2;
  logic [2:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR8;
  logic [131:0] zll_main_compute23_in;
  logic [130:0] zll_main_compute53_in;
  logic [7:0] zll_main_compute53_out;
  logic [130:0] zll_main_compute53_inR1;
  logic [7:0] zll_main_compute53_outR1;
  logic [130:0] zll_main_compute53_inR2;
  logic [7:0] zll_main_compute53_outR2;
  logic [130:0] zll_main_compute53_inR3;
  logic [7:0] zll_main_compute53_outR3;
  logic [130:0] zll_main_compute53_inR4;
  logic [7:0] zll_main_compute53_outR4;
  logic [130:0] zll_main_compute53_inR5;
  logic [7:0] zll_main_compute53_outR5;
  logic [130:0] zll_main_compute53_inR6;
  logic [7:0] zll_main_compute53_outR6;
  logic [130:0] zll_main_compute53_inR7;
  logic [7:0] zll_main_compute53_outR7;
  logic [63:0] resize_inR9;
  logic [2:0] resize_inR10;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR11;
  logic [2:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR13;
  assign resize_in = arg2;
  assign binop_in = {128'(resize_in[2:0]), 128'h3};
  assign resize_inR1 = arg2;
  assign binop_inR1 = {128'(resize_inR1[2:0]), 128'h3};
  assign zll_main_compute59_in = {arg2, arg0, arg1, binop_inR1[255:128] < binop_inR1[127:0]};
  assign zll_main_compute43_in = {zll_main_compute59_in[128:65], zll_main_compute59_in[64:1], 3'h0};
  ZLL_Main_compute43  inst (zll_main_compute43_in[130:67], zll_main_compute43_in[66:3], zll_main_compute43_in[2:0], zll_main_compute43_out);
  assign zll_main_compute43_inR1 = {zll_main_compute59_in[128:65], zll_main_compute59_in[64:1], 3'h1};
  ZLL_Main_compute43  instR1 (zll_main_compute43_inR1[130:67], zll_main_compute43_inR1[66:3], zll_main_compute43_inR1[2:0], zll_main_compute43_outR1);
  assign zll_main_compute43_inR2 = {zll_main_compute59_in[128:65], zll_main_compute59_in[64:1], 3'h2};
  ZLL_Main_compute43  instR2 (zll_main_compute43_inR2[130:67], zll_main_compute43_inR2[66:3], zll_main_compute43_inR2[2:0], zll_main_compute43_outR2);
  assign zll_main_compute43_inR3 = {zll_main_compute59_in[128:65], zll_main_compute59_in[64:1], 3'h3};
  ZLL_Main_compute43  instR3 (zll_main_compute43_inR3[130:67], zll_main_compute43_inR3[66:3], zll_main_compute43_inR3[2:0], zll_main_compute43_outR3);
  assign zll_main_compute43_inR4 = {zll_main_compute59_in[128:65], zll_main_compute59_in[64:1], 3'h4};
  ZLL_Main_compute43  instR4 (zll_main_compute43_inR4[130:67], zll_main_compute43_inR4[66:3], zll_main_compute43_inR4[2:0], zll_main_compute43_outR4);
  assign zll_main_compute43_inR5 = {zll_main_compute59_in[128:65], zll_main_compute59_in[64:1], 3'h5};
  ZLL_Main_compute43  instR5 (zll_main_compute43_inR5[130:67], zll_main_compute43_inR5[66:3], zll_main_compute43_inR5[2:0], zll_main_compute43_outR5);
  assign zll_main_compute43_inR6 = {zll_main_compute59_in[128:65], zll_main_compute59_in[64:1], 3'h6};
  ZLL_Main_compute43  instR6 (zll_main_compute43_inR6[130:67], zll_main_compute43_inR6[66:3], zll_main_compute43_inR6[2:0], zll_main_compute43_outR6);
  assign zll_main_compute43_inR7 = {zll_main_compute59_in[128:65], zll_main_compute59_in[64:1], 3'h7};
  ZLL_Main_compute43  instR7 (zll_main_compute43_inR7[130:67], zll_main_compute43_inR7[66:3], zll_main_compute43_inR7[2:0], zll_main_compute43_outR7);
  assign resize_inR2 = {zll_main_compute43_out, zll_main_compute43_outR1, zll_main_compute43_outR2, zll_main_compute43_outR3, zll_main_compute43_outR4, zll_main_compute43_outR5, zll_main_compute43_outR6, zll_main_compute43_outR7};
  assign resize_inR3 = zll_main_compute59_in[131:129];
  assign binop_inR2 = {128'(resize_inR3[2:0]), 128'h3};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h8};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[2:0];
  assign binop_inR4 = {128'(resize_inR5[2:0]), 128'h2};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h8};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR6 = {128'h8, 128'(resize_inR7[2:0])};
  assign binop_inR7 = {binop_inR6[255:128] - binop_inR6[127:0], 128'h1};
  assign binop_inR8 = {binop_inR7[255:128] - binop_inR7[127:0], 128'h8};
  assign binop_inR9 = {128'(resize_inR2[63:0]), binop_inR8[255:128] * binop_inR8[127:0]};
  assign resize_inR8 = binop_inR9[255:128] >> binop_inR9[127:0];
  assign zll_main_compute23_in = {arg2, arg0, arg1, binop_in[255:128] < binop_in[127:0]};
  assign zll_main_compute53_in = {zll_main_compute23_in[128:65], zll_main_compute23_in[64:1], 3'h0};
  ZLL_Main_compute53  instR8 (zll_main_compute53_in[130:67], zll_main_compute53_in[66:3], zll_main_compute53_in[2:0], zll_main_compute53_out);
  assign zll_main_compute53_inR1 = {zll_main_compute23_in[128:65], zll_main_compute23_in[64:1], 3'h1};
  ZLL_Main_compute53  instR9 (zll_main_compute53_inR1[130:67], zll_main_compute53_inR1[66:3], zll_main_compute53_inR1[2:0], zll_main_compute53_outR1);
  assign zll_main_compute53_inR2 = {zll_main_compute23_in[128:65], zll_main_compute23_in[64:1], 3'h2};
  ZLL_Main_compute53  instR10 (zll_main_compute53_inR2[130:67], zll_main_compute53_inR2[66:3], zll_main_compute53_inR2[2:0], zll_main_compute53_outR2);
  assign zll_main_compute53_inR3 = {zll_main_compute23_in[128:65], zll_main_compute23_in[64:1], 3'h3};
  ZLL_Main_compute53  instR11 (zll_main_compute53_inR3[130:67], zll_main_compute53_inR3[66:3], zll_main_compute53_inR3[2:0], zll_main_compute53_outR3);
  assign zll_main_compute53_inR4 = {zll_main_compute23_in[128:65], zll_main_compute23_in[64:1], 3'h4};
  ZLL_Main_compute53  instR12 (zll_main_compute53_inR4[130:67], zll_main_compute53_inR4[66:3], zll_main_compute53_inR4[2:0], zll_main_compute53_outR4);
  assign zll_main_compute53_inR5 = {zll_main_compute23_in[128:65], zll_main_compute23_in[64:1], 3'h5};
  ZLL_Main_compute53  instR13 (zll_main_compute53_inR5[130:67], zll_main_compute53_inR5[66:3], zll_main_compute53_inR5[2:0], zll_main_compute53_outR5);
  assign zll_main_compute53_inR6 = {zll_main_compute23_in[128:65], zll_main_compute23_in[64:1], 3'h6};
  ZLL_Main_compute53  instR14 (zll_main_compute53_inR6[130:67], zll_main_compute53_inR6[66:3], zll_main_compute53_inR6[2:0], zll_main_compute53_outR6);
  assign zll_main_compute53_inR7 = {zll_main_compute23_in[128:65], zll_main_compute23_in[64:1], 3'h7};
  ZLL_Main_compute53  instR15 (zll_main_compute53_inR7[130:67], zll_main_compute53_inR7[66:3], zll_main_compute53_inR7[2:0], zll_main_compute53_outR7);
  assign resize_inR9 = {zll_main_compute53_out, zll_main_compute53_outR1, zll_main_compute53_outR2, zll_main_compute53_outR3, zll_main_compute53_outR4, zll_main_compute53_outR5, zll_main_compute53_outR6, zll_main_compute53_outR7};
  assign resize_inR10 = zll_main_compute23_in[131:129];
  assign binop_inR10 = {128'(resize_inR10[2:0]), 128'h2};
  assign binop_inR11 = {binop_inR10[255:128] * binop_inR10[127:0], 128'h8};
  assign resize_inR11 = binop_inR11[255:128] % binop_inR11[127:0];
  assign resize_inR12 = resize_inR11[2:0];
  assign binop_inR12 = {128'h8, 128'(resize_inR12[2:0])};
  assign binop_inR13 = {binop_inR12[255:128] - binop_inR12[127:0], 128'h1};
  assign binop_inR14 = {binop_inR13[255:128] - binop_inR13[127:0], 128'h8};
  assign binop_inR15 = {128'(resize_inR9[63:0]), binop_inR14[255:128] * binop_inR14[127:0]};
  assign resize_inR13 = binop_inR15[255:128] >> binop_inR15[127:0];
  assign res = (zll_main_compute23_in[0] == 1'h1) ? resize_inR13[7:0] : resize_inR8[7:0];
endmodule

module ZLL_Main_compute34 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [127:0] resize_inR1;
  logic [0:0] msbit_in;
  logic [0:0] rewire_prelude_not_in;
  logic [0:0] rewire_prelude_not_out;
  logic [2:0] resize_inR2;
  logic [127:0] resize_inR3;
  logic [0:0] msbit_inR1;
  logic [0:0] rewire_prelude_not_inR1;
  logic [0:0] rewire_prelude_not_outR1;
  logic [131:0] zll_main_compute10_in;
  logic [130:0] zll_main_compute32_in;
  logic [7:0] zll_main_compute32_out;
  logic [130:0] zll_main_compute32_inR1;
  logic [7:0] zll_main_compute32_outR1;
  logic [130:0] zll_main_compute32_inR2;
  logic [7:0] zll_main_compute32_outR2;
  logic [130:0] zll_main_compute32_inR3;
  logic [7:0] zll_main_compute32_outR3;
  logic [130:0] zll_main_compute32_inR4;
  logic [7:0] zll_main_compute32_outR4;
  logic [130:0] zll_main_compute32_inR5;
  logic [7:0] zll_main_compute32_outR5;
  logic [130:0] zll_main_compute32_inR6;
  logic [7:0] zll_main_compute32_outR6;
  logic [130:0] zll_main_compute32_inR7;
  logic [7:0] zll_main_compute32_outR7;
  logic [63:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR8;
  logic [2:0] resize_inR9;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR10;
  logic [2:0] resize_inR11;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [127:0] resize_inR12;
  logic [131:0] zll_main_compute20_in;
  logic [130:0] zll_main_compute36_in;
  logic [7:0] zll_main_compute36_out;
  logic [130:0] zll_main_compute36_inR1;
  logic [7:0] zll_main_compute36_outR1;
  logic [130:0] zll_main_compute36_inR2;
  logic [7:0] zll_main_compute36_outR2;
  logic [130:0] zll_main_compute36_inR3;
  logic [7:0] zll_main_compute36_outR3;
  logic [130:0] zll_main_compute36_inR4;
  logic [7:0] zll_main_compute36_outR4;
  logic [130:0] zll_main_compute36_inR5;
  logic [7:0] zll_main_compute36_outR5;
  logic [130:0] zll_main_compute36_inR6;
  logic [7:0] zll_main_compute36_outR6;
  logic [130:0] zll_main_compute36_inR7;
  logic [7:0] zll_main_compute36_outR7;
  logic [63:0] resize_inR13;
  logic [2:0] resize_inR14;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR15;
  logic [2:0] resize_inR16;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [127:0] resize_inR17;
  logic [2:0] resize_inR18;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [255:0] binop_inR16;
  logic [255:0] binop_inR17;
  logic [127:0] resize_inR19;
  assign resize_in = arg2;
  assign resize_inR1 = 128'(resize_in[2:0]);
  assign msbit_in = resize_inR1[0];
  assign rewire_prelude_not_in = msbit_in[0];
  ReWire_Prelude_not  inst (rewire_prelude_not_in[0], rewire_prelude_not_out);
  assign resize_inR2 = arg2;
  assign resize_inR3 = 128'(resize_inR2[2:0]);
  assign msbit_inR1 = resize_inR3[0];
  assign rewire_prelude_not_inR1 = msbit_inR1[0];
  ReWire_Prelude_not  instR1 (rewire_prelude_not_inR1[0], rewire_prelude_not_outR1);
  assign zll_main_compute10_in = {arg0, arg1, arg2, rewire_prelude_not_outR1};
  assign zll_main_compute32_in = {zll_main_compute10_in[131:68], zll_main_compute10_in[67:4], 3'h0};
  ZLL_Main_compute32  instR2 (zll_main_compute32_in[130:67], zll_main_compute32_in[66:3], zll_main_compute32_in[2:0], zll_main_compute32_out);
  assign zll_main_compute32_inR1 = {zll_main_compute10_in[131:68], zll_main_compute10_in[67:4], 3'h1};
  ZLL_Main_compute32  instR3 (zll_main_compute32_inR1[130:67], zll_main_compute32_inR1[66:3], zll_main_compute32_inR1[2:0], zll_main_compute32_outR1);
  assign zll_main_compute32_inR2 = {zll_main_compute10_in[131:68], zll_main_compute10_in[67:4], 3'h2};
  ZLL_Main_compute32  instR4 (zll_main_compute32_inR2[130:67], zll_main_compute32_inR2[66:3], zll_main_compute32_inR2[2:0], zll_main_compute32_outR2);
  assign zll_main_compute32_inR3 = {zll_main_compute10_in[131:68], zll_main_compute10_in[67:4], 3'h3};
  ZLL_Main_compute32  instR5 (zll_main_compute32_inR3[130:67], zll_main_compute32_inR3[66:3], zll_main_compute32_inR3[2:0], zll_main_compute32_outR3);
  assign zll_main_compute32_inR4 = {zll_main_compute10_in[131:68], zll_main_compute10_in[67:4], 3'h4};
  ZLL_Main_compute32  instR6 (zll_main_compute32_inR4[130:67], zll_main_compute32_inR4[66:3], zll_main_compute32_inR4[2:0], zll_main_compute32_outR4);
  assign zll_main_compute32_inR5 = {zll_main_compute10_in[131:68], zll_main_compute10_in[67:4], 3'h5};
  ZLL_Main_compute32  instR7 (zll_main_compute32_inR5[130:67], zll_main_compute32_inR5[66:3], zll_main_compute32_inR5[2:0], zll_main_compute32_outR5);
  assign zll_main_compute32_inR6 = {zll_main_compute10_in[131:68], zll_main_compute10_in[67:4], 3'h6};
  ZLL_Main_compute32  instR8 (zll_main_compute32_inR6[130:67], zll_main_compute32_inR6[66:3], zll_main_compute32_inR6[2:0], zll_main_compute32_outR6);
  assign zll_main_compute32_inR7 = {zll_main_compute10_in[131:68], zll_main_compute10_in[67:4], 3'h7};
  ZLL_Main_compute32  instR9 (zll_main_compute32_inR7[130:67], zll_main_compute32_inR7[66:3], zll_main_compute32_inR7[2:0], zll_main_compute32_outR7);
  assign resize_inR4 = {zll_main_compute32_out, zll_main_compute32_outR1, zll_main_compute32_outR2, zll_main_compute32_outR3, zll_main_compute32_outR4, zll_main_compute32_outR5, zll_main_compute32_outR6, zll_main_compute32_outR7};
  assign resize_inR5 = zll_main_compute10_in[3:1];
  assign binop_in = {128'(resize_inR5[2:0]), 128'h1};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h8};
  assign resize_inR6 = binop_inR1[255:128] % binop_inR1[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR2 = {128'h3, 128'(resize_inR7[2:0])};
  assign binop_inR3 = {binop_inR2[255:128] + binop_inR2[127:0], 128'h8};
  assign resize_inR8 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR9 = resize_inR8[2:0];
  assign binop_inR4 = {128'(resize_inR9[2:0]), 128'h2};
  assign binop_inR5 = {binop_inR4[255:128] / binop_inR4[127:0], 128'h8};
  assign resize_inR10 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR11 = resize_inR10[2:0];
  assign binop_inR6 = {128'h8, 128'(resize_inR11[2:0])};
  assign binop_inR7 = {binop_inR6[255:128] - binop_inR6[127:0], 128'h1};
  assign binop_inR8 = {binop_inR7[255:128] - binop_inR7[127:0], 128'h8};
  assign binop_inR9 = {128'(resize_inR4[63:0]), binop_inR8[255:128] * binop_inR8[127:0]};
  assign resize_inR12 = binop_inR9[255:128] >> binop_inR9[127:0];
  assign zll_main_compute20_in = {arg0, arg1, arg2, rewire_prelude_not_out};
  assign zll_main_compute36_in = {zll_main_compute20_in[131:68], zll_main_compute20_in[67:4], 3'h0};
  ZLL_Main_compute36  instR10 (zll_main_compute36_in[130:67], zll_main_compute36_in[66:3], zll_main_compute36_in[2:0], zll_main_compute36_out);
  assign zll_main_compute36_inR1 = {zll_main_compute20_in[131:68], zll_main_compute20_in[67:4], 3'h1};
  ZLL_Main_compute36  instR11 (zll_main_compute36_inR1[130:67], zll_main_compute36_inR1[66:3], zll_main_compute36_inR1[2:0], zll_main_compute36_outR1);
  assign zll_main_compute36_inR2 = {zll_main_compute20_in[131:68], zll_main_compute20_in[67:4], 3'h2};
  ZLL_Main_compute36  instR12 (zll_main_compute36_inR2[130:67], zll_main_compute36_inR2[66:3], zll_main_compute36_inR2[2:0], zll_main_compute36_outR2);
  assign zll_main_compute36_inR3 = {zll_main_compute20_in[131:68], zll_main_compute20_in[67:4], 3'h3};
  ZLL_Main_compute36  instR13 (zll_main_compute36_inR3[130:67], zll_main_compute36_inR3[66:3], zll_main_compute36_inR3[2:0], zll_main_compute36_outR3);
  assign zll_main_compute36_inR4 = {zll_main_compute20_in[131:68], zll_main_compute20_in[67:4], 3'h4};
  ZLL_Main_compute36  instR14 (zll_main_compute36_inR4[130:67], zll_main_compute36_inR4[66:3], zll_main_compute36_inR4[2:0], zll_main_compute36_outR4);
  assign zll_main_compute36_inR5 = {zll_main_compute20_in[131:68], zll_main_compute20_in[67:4], 3'h5};
  ZLL_Main_compute36  instR15 (zll_main_compute36_inR5[130:67], zll_main_compute36_inR5[66:3], zll_main_compute36_inR5[2:0], zll_main_compute36_outR5);
  assign zll_main_compute36_inR6 = {zll_main_compute20_in[131:68], zll_main_compute20_in[67:4], 3'h6};
  ZLL_Main_compute36  instR16 (zll_main_compute36_inR6[130:67], zll_main_compute36_inR6[66:3], zll_main_compute36_inR6[2:0], zll_main_compute36_outR6);
  assign zll_main_compute36_inR7 = {zll_main_compute20_in[131:68], zll_main_compute20_in[67:4], 3'h7};
  ZLL_Main_compute36  instR17 (zll_main_compute36_inR7[130:67], zll_main_compute36_inR7[66:3], zll_main_compute36_inR7[2:0], zll_main_compute36_outR7);
  assign resize_inR13 = {zll_main_compute36_out, zll_main_compute36_outR1, zll_main_compute36_outR2, zll_main_compute36_outR3, zll_main_compute36_outR4, zll_main_compute36_outR5, zll_main_compute36_outR6, zll_main_compute36_outR7};
  assign resize_inR14 = zll_main_compute20_in[3:1];
  assign binop_inR10 = {128'h3, 128'(resize_inR14[2:0])};
  assign binop_inR11 = {binop_inR10[255:128] + binop_inR10[127:0], 128'h8};
  assign resize_inR15 = binop_inR11[255:128] % binop_inR11[127:0];
  assign resize_inR16 = resize_inR15[2:0];
  assign binop_inR12 = {128'(resize_inR16[2:0]), 128'h2};
  assign binop_inR13 = {binop_inR12[255:128] / binop_inR12[127:0], 128'h8};
  assign resize_inR17 = binop_inR13[255:128] % binop_inR13[127:0];
  assign resize_inR18 = resize_inR17[2:0];
  assign binop_inR14 = {128'h8, 128'(resize_inR18[2:0])};
  assign binop_inR15 = {binop_inR14[255:128] - binop_inR14[127:0], 128'h1};
  assign binop_inR16 = {binop_inR15[255:128] - binop_inR15[127:0], 128'h8};
  assign binop_inR17 = {128'(resize_inR13[63:0]), binop_inR16[255:128] * binop_inR16[127:0]};
  assign resize_inR19 = binop_inR17[255:128] >> binop_inR17[127:0];
  assign res = (zll_main_compute20_in[0] == 1'h1) ? resize_inR19[7:0] : resize_inR12[7:0];
endmodule

module ZLL_Main_compute32 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resize_in;
  logic [255:0] binop_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_inR1;
  logic [131:0] zll_main_compute85_in;
  logic [130:0] zll_main_compute43_in;
  logic [7:0] zll_main_compute43_out;
  logic [130:0] zll_main_compute43_inR1;
  logic [7:0] zll_main_compute43_outR1;
  logic [130:0] zll_main_compute43_inR2;
  logic [7:0] zll_main_compute43_outR2;
  logic [130:0] zll_main_compute43_inR3;
  logic [7:0] zll_main_compute43_outR3;
  logic [130:0] zll_main_compute43_inR4;
  logic [7:0] zll_main_compute43_outR4;
  logic [130:0] zll_main_compute43_inR5;
  logic [7:0] zll_main_compute43_outR5;
  logic [130:0] zll_main_compute43_inR6;
  logic [7:0] zll_main_compute43_outR6;
  logic [130:0] zll_main_compute43_inR7;
  logic [7:0] zll_main_compute43_outR7;
  logic [63:0] resize_inR2;
  logic [2:0] resize_inR3;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR4;
  logic [2:0] resize_inR5;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [127:0] resize_inR6;
  logic [2:0] resize_inR7;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR8;
  logic [2:0] resize_inR9;
  logic [255:0] binop_inR8;
  logic [255:0] binop_inR9;
  logic [255:0] binop_inR10;
  logic [255:0] binop_inR11;
  logic [127:0] resize_inR10;
  logic [131:0] zll_main_compute79_in;
  logic [130:0] zll_main_compute53_in;
  logic [7:0] zll_main_compute53_out;
  logic [130:0] zll_main_compute53_inR1;
  logic [7:0] zll_main_compute53_outR1;
  logic [130:0] zll_main_compute53_inR2;
  logic [7:0] zll_main_compute53_outR2;
  logic [130:0] zll_main_compute53_inR3;
  logic [7:0] zll_main_compute53_outR3;
  logic [130:0] zll_main_compute53_inR4;
  logic [7:0] zll_main_compute53_outR4;
  logic [130:0] zll_main_compute53_inR5;
  logic [7:0] zll_main_compute53_outR5;
  logic [130:0] zll_main_compute53_inR6;
  logic [7:0] zll_main_compute53_outR6;
  logic [130:0] zll_main_compute53_inR7;
  logic [7:0] zll_main_compute53_outR7;
  logic [63:0] resize_inR11;
  logic [2:0] resize_inR12;
  logic [255:0] binop_inR12;
  logic [255:0] binop_inR13;
  logic [127:0] resize_inR13;
  logic [2:0] resize_inR14;
  logic [255:0] binop_inR14;
  logic [255:0] binop_inR15;
  logic [127:0] resize_inR15;
  logic [2:0] resize_inR16;
  logic [255:0] binop_inR16;
  logic [255:0] binop_inR17;
  logic [255:0] binop_inR18;
  logic [255:0] binop_inR19;
  logic [127:0] resize_inR17;
  assign resize_in = arg2;
  assign binop_in = {128'(resize_in[2:0]), 128'h3};
  assign resize_inR1 = arg2;
  assign binop_inR1 = {128'(resize_inR1[2:0]), 128'h3};
  assign zll_main_compute85_in = {arg2, arg0, arg1, binop_inR1[255:128] < binop_inR1[127:0]};
  assign zll_main_compute43_in = {zll_main_compute85_in[128:65], zll_main_compute85_in[64:1], 3'h0};
  ZLL_Main_compute43  inst (zll_main_compute43_in[130:67], zll_main_compute43_in[66:3], zll_main_compute43_in[2:0], zll_main_compute43_out);
  assign zll_main_compute43_inR1 = {zll_main_compute85_in[128:65], zll_main_compute85_in[64:1], 3'h1};
  ZLL_Main_compute43  instR1 (zll_main_compute43_inR1[130:67], zll_main_compute43_inR1[66:3], zll_main_compute43_inR1[2:0], zll_main_compute43_outR1);
  assign zll_main_compute43_inR2 = {zll_main_compute85_in[128:65], zll_main_compute85_in[64:1], 3'h2};
  ZLL_Main_compute43  instR2 (zll_main_compute43_inR2[130:67], zll_main_compute43_inR2[66:3], zll_main_compute43_inR2[2:0], zll_main_compute43_outR2);
  assign zll_main_compute43_inR3 = {zll_main_compute85_in[128:65], zll_main_compute85_in[64:1], 3'h3};
  ZLL_Main_compute43  instR3 (zll_main_compute43_inR3[130:67], zll_main_compute43_inR3[66:3], zll_main_compute43_inR3[2:0], zll_main_compute43_outR3);
  assign zll_main_compute43_inR4 = {zll_main_compute85_in[128:65], zll_main_compute85_in[64:1], 3'h4};
  ZLL_Main_compute43  instR4 (zll_main_compute43_inR4[130:67], zll_main_compute43_inR4[66:3], zll_main_compute43_inR4[2:0], zll_main_compute43_outR4);
  assign zll_main_compute43_inR5 = {zll_main_compute85_in[128:65], zll_main_compute85_in[64:1], 3'h5};
  ZLL_Main_compute43  instR5 (zll_main_compute43_inR5[130:67], zll_main_compute43_inR5[66:3], zll_main_compute43_inR5[2:0], zll_main_compute43_outR5);
  assign zll_main_compute43_inR6 = {zll_main_compute85_in[128:65], zll_main_compute85_in[64:1], 3'h6};
  ZLL_Main_compute43  instR6 (zll_main_compute43_inR6[130:67], zll_main_compute43_inR6[66:3], zll_main_compute43_inR6[2:0], zll_main_compute43_outR6);
  assign zll_main_compute43_inR7 = {zll_main_compute85_in[128:65], zll_main_compute85_in[64:1], 3'h7};
  ZLL_Main_compute43  instR7 (zll_main_compute43_inR7[130:67], zll_main_compute43_inR7[66:3], zll_main_compute43_inR7[2:0], zll_main_compute43_outR7);
  assign resize_inR2 = {zll_main_compute43_out, zll_main_compute43_outR1, zll_main_compute43_outR2, zll_main_compute43_outR3, zll_main_compute43_outR4, zll_main_compute43_outR5, zll_main_compute43_outR6, zll_main_compute43_outR7};
  assign resize_inR3 = zll_main_compute85_in[131:129];
  assign binop_inR2 = {128'(resize_inR3[2:0]), 128'h3};
  assign binop_inR3 = {binop_inR2[255:128] - binop_inR2[127:0], 128'h8};
  assign resize_inR4 = binop_inR3[255:128] % binop_inR3[127:0];
  assign resize_inR5 = resize_inR4[2:0];
  assign binop_inR4 = {128'(resize_inR5[2:0]), 128'h2};
  assign binop_inR5 = {binop_inR4[255:128] * binop_inR4[127:0], 128'h8};
  assign resize_inR6 = binop_inR5[255:128] % binop_inR5[127:0];
  assign resize_inR7 = resize_inR6[2:0];
  assign binop_inR6 = {128'(resize_inR7[2:0]), 128'h1};
  assign binop_inR7 = {binop_inR6[255:128] + binop_inR6[127:0], 128'h8};
  assign resize_inR8 = binop_inR7[255:128] % binop_inR7[127:0];
  assign resize_inR9 = resize_inR8[2:0];
  assign binop_inR8 = {128'h8, 128'(resize_inR9[2:0])};
  assign binop_inR9 = {binop_inR8[255:128] - binop_inR8[127:0], 128'h1};
  assign binop_inR10 = {binop_inR9[255:128] - binop_inR9[127:0], 128'h8};
  assign binop_inR11 = {128'(resize_inR2[63:0]), binop_inR10[255:128] * binop_inR10[127:0]};
  assign resize_inR10 = binop_inR11[255:128] >> binop_inR11[127:0];
  assign zll_main_compute79_in = {arg2, arg0, arg1, binop_in[255:128] < binop_in[127:0]};
  assign zll_main_compute53_in = {zll_main_compute79_in[128:65], zll_main_compute79_in[64:1], 3'h0};
  ZLL_Main_compute53  instR8 (zll_main_compute53_in[130:67], zll_main_compute53_in[66:3], zll_main_compute53_in[2:0], zll_main_compute53_out);
  assign zll_main_compute53_inR1 = {zll_main_compute79_in[128:65], zll_main_compute79_in[64:1], 3'h1};
  ZLL_Main_compute53  instR9 (zll_main_compute53_inR1[130:67], zll_main_compute53_inR1[66:3], zll_main_compute53_inR1[2:0], zll_main_compute53_outR1);
  assign zll_main_compute53_inR2 = {zll_main_compute79_in[128:65], zll_main_compute79_in[64:1], 3'h2};
  ZLL_Main_compute53  instR10 (zll_main_compute53_inR2[130:67], zll_main_compute53_inR2[66:3], zll_main_compute53_inR2[2:0], zll_main_compute53_outR2);
  assign zll_main_compute53_inR3 = {zll_main_compute79_in[128:65], zll_main_compute79_in[64:1], 3'h3};
  ZLL_Main_compute53  instR11 (zll_main_compute53_inR3[130:67], zll_main_compute53_inR3[66:3], zll_main_compute53_inR3[2:0], zll_main_compute53_outR3);
  assign zll_main_compute53_inR4 = {zll_main_compute79_in[128:65], zll_main_compute79_in[64:1], 3'h4};
  ZLL_Main_compute53  instR12 (zll_main_compute53_inR4[130:67], zll_main_compute53_inR4[66:3], zll_main_compute53_inR4[2:0], zll_main_compute53_outR4);
  assign zll_main_compute53_inR5 = {zll_main_compute79_in[128:65], zll_main_compute79_in[64:1], 3'h5};
  ZLL_Main_compute53  instR13 (zll_main_compute53_inR5[130:67], zll_main_compute53_inR5[66:3], zll_main_compute53_inR5[2:0], zll_main_compute53_outR5);
  assign zll_main_compute53_inR6 = {zll_main_compute79_in[128:65], zll_main_compute79_in[64:1], 3'h6};
  ZLL_Main_compute53  instR14 (zll_main_compute53_inR6[130:67], zll_main_compute53_inR6[66:3], zll_main_compute53_inR6[2:0], zll_main_compute53_outR6);
  assign zll_main_compute53_inR7 = {zll_main_compute79_in[128:65], zll_main_compute79_in[64:1], 3'h7};
  ZLL_Main_compute53  instR15 (zll_main_compute53_inR7[130:67], zll_main_compute53_inR7[66:3], zll_main_compute53_inR7[2:0], zll_main_compute53_outR7);
  assign resize_inR11 = {zll_main_compute53_out, zll_main_compute53_outR1, zll_main_compute53_outR2, zll_main_compute53_outR3, zll_main_compute53_outR4, zll_main_compute53_outR5, zll_main_compute53_outR6, zll_main_compute53_outR7};
  assign resize_inR12 = zll_main_compute79_in[131:129];
  assign binop_inR12 = {128'(resize_inR12[2:0]), 128'h2};
  assign binop_inR13 = {binop_inR12[255:128] * binop_inR12[127:0], 128'h8};
  assign resize_inR13 = binop_inR13[255:128] % binop_inR13[127:0];
  assign resize_inR14 = resize_inR13[2:0];
  assign binop_inR14 = {128'(resize_inR14[2:0]), 128'h1};
  assign binop_inR15 = {binop_inR14[255:128] + binop_inR14[127:0], 128'h8};
  assign resize_inR15 = binop_inR15[255:128] % binop_inR15[127:0];
  assign resize_inR16 = resize_inR15[2:0];
  assign binop_inR16 = {128'h8, 128'(resize_inR16[2:0])};
  assign binop_inR17 = {binop_inR16[255:128] - binop_inR16[127:0], 128'h1};
  assign binop_inR18 = {binop_inR17[255:128] - binop_inR17[127:0], 128'h8};
  assign binop_inR19 = {128'(resize_inR11[63:0]), binop_inR18[255:128] * binop_inR18[127:0]};
  assign resize_inR17 = binop_inR19[255:128] >> binop_inR19[127:0];
  assign res = (zll_main_compute79_in[0] == 1'h1) ? resize_inR17[7:0] : resize_inR10[7:0];
endmodule