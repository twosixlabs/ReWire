module top_level ();
  logic [0:0] __continue;
endmodule