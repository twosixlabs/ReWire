module top_level (input logic [63:0] __in0,
  input logic [63:0] __in1,
  output logic [63:0] __out0,
  output logic [63:0] __out1);
  logic [127:0] zll_main_loop3_in;
  logic [127:0] zll_main_compute66_in;
  logic [127:0] zll_main_compute191_in;
  logic [127:0] zll_main_compute270_in;
  logic [127:0] zll_main_compute67_in;
  logic [127:0] zll_main_compute83_in;
  logic [130:0] zll_main_compute307_in;
  logic [133:0] zll_main_compute102_in;
  logic [5:0] zll_main_compute428_in;
  logic [2:0] zll_main_compute428_out;
  logic [136:0] zll_main_compute267_in;
  logic [70:0] zll_main_compute418_in;
  logic [6:0] zll_main_compute354_in;
  logic [2:0] zll_main_compute354_out;
  logic [3:0] id_in;
  logic [133:0] zll_main_compute57_in;
  logic [136:0] zll_main_compute259_in;
  logic [7:0] zll_main_compute259_out;
  logic [136:0] zll_main_compute259_inR1;
  logic [7:0] zll_main_compute259_outR1;
  logic [136:0] zll_main_compute259_inR2;
  logic [7:0] zll_main_compute259_outR2;
  logic [136:0] zll_main_compute259_inR3;
  logic [7:0] zll_main_compute259_outR3;
  logic [136:0] zll_main_compute259_inR4;
  logic [7:0] zll_main_compute259_outR4;
  logic [136:0] zll_main_compute259_inR5;
  logic [7:0] zll_main_compute259_outR5;
  logic [136:0] zll_main_compute259_inR6;
  logic [7:0] zll_main_compute259_outR6;
  logic [136:0] zll_main_compute259_inR7;
  logic [7:0] zll_main_compute259_outR7;
  logic [127:0] zll_main_compute124_in;
  logic [127:0] zll_main_compute190_in;
  logic [127:0] zll_main_compute375_in;
  logic [127:0] zll_main_compute31_in;
  logic [130:0] zll_main_compute148_in;
  logic [133:0] zll_main_compute353_in;
  logic [5:0] zll_main_compute428_inR1;
  logic [2:0] zll_main_compute428_outR1;
  logic [136:0] zll_main_compute70_in;
  logic [70:0] zll_main_compute383_in;
  logic [2:0] zll_main_compute383_out;
  logic [136:0] zll_main_compute275_in;
  logic [139:0] zll_main_compute119_in;
  logic [7:0] zll_main_compute119_out;
  logic [139:0] zll_main_compute119_inR1;
  logic [7:0] zll_main_compute119_outR1;
  logic [139:0] zll_main_compute119_inR2;
  logic [7:0] zll_main_compute119_outR2;
  logic [139:0] zll_main_compute119_inR3;
  logic [7:0] zll_main_compute119_outR3;
  logic [139:0] zll_main_compute119_inR4;
  logic [7:0] zll_main_compute119_outR4;
  logic [139:0] zll_main_compute119_inR5;
  logic [7:0] zll_main_compute119_outR5;
  logic [139:0] zll_main_compute119_inR6;
  logic [7:0] zll_main_compute119_outR6;
  logic [139:0] zll_main_compute119_inR7;
  logic [7:0] zll_main_compute119_outR7;
  logic [127:0] zll_main_compute329_in;
  logic [127:0] zll_main_compute232_in;
  logic [127:0] zll_main_compute365_in;
  logic [127:0] zll_main_compute254_in;
  logic [127:0] zll_main_compute80_in;
  logic [130:0] zll_main_compute183_in;
  logic [130:0] zll_main_compute422_in;
  logic [133:0] zll_main_compute417_in;
  logic [5:0] zll_main_compute428_inR2;
  logic [2:0] zll_main_compute428_outR2;
  logic [136:0] zll_main_compute348_in;
  logic [70:0] zll_main_compute6_in;
  logic [6:0] zll_main_compute354_inR1;
  logic [2:0] zll_main_compute354_outR1;
  logic [3:0] id_inR1;
  logic [133:0] zll_main_compute118_in;
  logic [136:0] zll_main_compute221_in;
  logic [7:0] zll_main_compute221_out;
  logic [136:0] zll_main_compute221_inR1;
  logic [7:0] zll_main_compute221_outR1;
  logic [136:0] zll_main_compute221_inR2;
  logic [7:0] zll_main_compute221_outR2;
  logic [136:0] zll_main_compute221_inR3;
  logic [7:0] zll_main_compute221_outR3;
  logic [136:0] zll_main_compute221_inR4;
  logic [7:0] zll_main_compute221_outR4;
  logic [136:0] zll_main_compute221_inR5;
  logic [7:0] zll_main_compute221_outR5;
  logic [136:0] zll_main_compute221_inR6;
  logic [7:0] zll_main_compute221_outR6;
  logic [136:0] zll_main_compute221_inR7;
  logic [7:0] zll_main_compute221_outR7;
  logic [127:0] zll_main_compute180_in;
  logic [127:0] zll_main_compute20_in;
  logic [127:0] zll_main_compute441_in;
  logic [127:0] zll_main_compute437_in;
  logic [130:0] zll_main_compute324_in;
  logic [130:0] zll_main_compute396_in;
  logic [133:0] zll_main_compute398_in;
  logic [5:0] zll_main_compute428_inR3;
  logic [2:0] zll_main_compute428_outR3;
  logic [136:0] zll_main_compute407_in;
  logic [70:0] zll_main_compute351_in;
  logic [6:0] zll_main_compute321_in;
  logic [2:0] zll_main_compute321_out;
  logic [3:0] id_inR2;
  logic [136:0] zll_main_compute16_in;
  logic [139:0] zll_main_compute28_in;
  logic [7:0] zll_main_compute28_out;
  logic [139:0] zll_main_compute28_inR1;
  logic [7:0] zll_main_compute28_outR1;
  logic [139:0] zll_main_compute28_inR2;
  logic [7:0] zll_main_compute28_outR2;
  logic [139:0] zll_main_compute28_inR3;
  logic [7:0] zll_main_compute28_outR3;
  logic [139:0] zll_main_compute28_inR4;
  logic [7:0] zll_main_compute28_outR4;
  logic [139:0] zll_main_compute28_inR5;
  logic [7:0] zll_main_compute28_outR5;
  logic [139:0] zll_main_compute28_inR6;
  logic [7:0] zll_main_compute28_outR6;
  logic [139:0] zll_main_compute28_inR7;
  logic [7:0] zll_main_compute28_outR7;
  logic [127:0] zll_main_compute97_in;
  logic [127:0] zll_main_compute357_in;
  logic [127:0] zll_main_compute293_in;
  logic [127:0] zll_main_compute371_in;
  logic [127:0] zll_main_compute160_in;
  logic [127:0] zll_main_compute279_in;
  logic [130:0] zll_main_compute178_in;
  logic [133:0] zll_main_compute261_in;
  logic [136:0] zll_main_compute198_in;
  logic [7:0] zll_main_compute198_out;
  logic [136:0] zll_main_compute198_inR1;
  logic [7:0] zll_main_compute198_outR1;
  logic [136:0] zll_main_compute198_inR2;
  logic [7:0] zll_main_compute198_outR2;
  logic [136:0] zll_main_compute198_inR3;
  logic [7:0] zll_main_compute198_outR3;
  logic [136:0] zll_main_compute198_inR4;
  logic [7:0] zll_main_compute198_outR4;
  logic [136:0] zll_main_compute198_inR5;
  logic [7:0] zll_main_compute198_outR5;
  logic [136:0] zll_main_compute198_inR6;
  logic [7:0] zll_main_compute198_outR6;
  logic [136:0] zll_main_compute198_inR7;
  logic [7:0] zll_main_compute198_outR7;
  logic [127:0] zll_main_compute286_in;
  logic [127:0] zll_main_compute127_in;
  logic [127:0] zll_main_compute399_in;
  logic [130:0] zll_main_compute243_in;
  logic [133:0] zll_main_compute55_in;
  logic [5:0] zll_main_compute428_inR4;
  logic [2:0] zll_main_compute428_outR4;
  logic [136:0] zll_main_compute96_in;
  logic [70:0] zll_main_compute383_inR1;
  logic [2:0] zll_main_compute383_outR1;
  logic [136:0] zll_main_compute406_in;
  logic [139:0] zll_main_compute141_in;
  logic [7:0] zll_main_compute141_out;
  logic [139:0] zll_main_compute141_inR1;
  logic [7:0] zll_main_compute141_outR1;
  logic [139:0] zll_main_compute141_inR2;
  logic [7:0] zll_main_compute141_outR2;
  logic [139:0] zll_main_compute141_inR3;
  logic [7:0] zll_main_compute141_outR3;
  logic [139:0] zll_main_compute141_inR4;
  logic [7:0] zll_main_compute141_outR4;
  logic [139:0] zll_main_compute141_inR5;
  logic [7:0] zll_main_compute141_outR5;
  logic [139:0] zll_main_compute141_inR6;
  logic [7:0] zll_main_compute141_outR6;
  logic [139:0] zll_main_compute141_inR7;
  logic [7:0] zll_main_compute141_outR7;
  logic [127:0] zll_main_compute442_in;
  logic [127:0] id_inR3;
  logic [128:0] zll_main_loop1_in;
  logic [128:0] zll_main_loop2_in;
  logic [0:0] __continue;
  assign zll_main_loop3_in = {__in0, __in1};
  assign zll_main_compute66_in = zll_main_loop3_in[127:0];
  assign zll_main_compute191_in = zll_main_compute66_in[127:0];
  assign zll_main_compute270_in = {zll_main_compute191_in[127:64], zll_main_compute191_in[63:0]};
  assign zll_main_compute67_in = {zll_main_compute270_in[127:64], zll_main_compute270_in[63:0]};
  assign zll_main_compute83_in = zll_main_compute67_in[127:0];
  assign zll_main_compute307_in = {zll_main_compute83_in[127:64], zll_main_compute83_in[63:0], 3'h1};
  assign zll_main_compute102_in = {zll_main_compute307_in[130:67], zll_main_compute307_in[66:3], zll_main_compute307_in[2:0], 3'h2};
  assign zll_main_compute428_in = {3'h7, zll_main_compute102_in[2:0]};
  ZLL_Main_compute428  inst (zll_main_compute428_in[5:3], zll_main_compute428_in[2:0], zll_main_compute428_out);
  assign zll_main_compute267_in = {zll_main_compute102_in[133:70], zll_main_compute102_in[69:6], zll_main_compute102_in[2:0], zll_main_compute102_in[5:3], zll_main_compute428_out};
  assign zll_main_compute418_in = {zll_main_compute267_in[136:73], zll_main_compute267_in[5:3], zll_main_compute267_in[2:0], 1'h0};
  assign zll_main_compute354_in = {zll_main_compute418_in[6:4], zll_main_compute418_in[3:1], 1'h0};
  ZLL_Main_compute354  instR1 (zll_main_compute354_in[6:4], zll_main_compute354_in[3:1], zll_main_compute354_in[0], zll_main_compute354_out);
  assign id_in = {zll_main_compute418_in[3:1], zll_main_compute418_in[0]};
  assign zll_main_compute57_in = {zll_main_compute267_in[136:73], zll_main_compute267_in[72:9], zll_main_compute267_in[8:6], (id_in[0] == 1'h1) ? id_in[3:1] : zll_main_compute354_out};
  assign zll_main_compute259_in = {zll_main_compute57_in[133:70], zll_main_compute57_in[69:6], zll_main_compute57_in[5:3], zll_main_compute57_in[2:0], 3'h0};
  ZLL_Main_compute259  instR2 (zll_main_compute259_in[136:73], zll_main_compute259_in[72:9], zll_main_compute259_in[8:6], zll_main_compute259_in[5:3], zll_main_compute259_in[2:0], zll_main_compute259_out);
  assign zll_main_compute259_inR1 = {zll_main_compute57_in[133:70], zll_main_compute57_in[69:6], zll_main_compute57_in[5:3], zll_main_compute57_in[2:0], 3'h1};
  ZLL_Main_compute259  instR3 (zll_main_compute259_inR1[136:73], zll_main_compute259_inR1[72:9], zll_main_compute259_inR1[8:6], zll_main_compute259_inR1[5:3], zll_main_compute259_inR1[2:0], zll_main_compute259_outR1);
  assign zll_main_compute259_inR2 = {zll_main_compute57_in[133:70], zll_main_compute57_in[69:6], zll_main_compute57_in[5:3], zll_main_compute57_in[2:0], 3'h2};
  ZLL_Main_compute259  instR4 (zll_main_compute259_inR2[136:73], zll_main_compute259_inR2[72:9], zll_main_compute259_inR2[8:6], zll_main_compute259_inR2[5:3], zll_main_compute259_inR2[2:0], zll_main_compute259_outR2);
  assign zll_main_compute259_inR3 = {zll_main_compute57_in[133:70], zll_main_compute57_in[69:6], zll_main_compute57_in[5:3], zll_main_compute57_in[2:0], 3'h3};
  ZLL_Main_compute259  instR5 (zll_main_compute259_inR3[136:73], zll_main_compute259_inR3[72:9], zll_main_compute259_inR3[8:6], zll_main_compute259_inR3[5:3], zll_main_compute259_inR3[2:0], zll_main_compute259_outR3);
  assign zll_main_compute259_inR4 = {zll_main_compute57_in[133:70], zll_main_compute57_in[69:6], zll_main_compute57_in[5:3], zll_main_compute57_in[2:0], 3'h4};
  ZLL_Main_compute259  instR6 (zll_main_compute259_inR4[136:73], zll_main_compute259_inR4[72:9], zll_main_compute259_inR4[8:6], zll_main_compute259_inR4[5:3], zll_main_compute259_inR4[2:0], zll_main_compute259_outR4);
  assign zll_main_compute259_inR5 = {zll_main_compute57_in[133:70], zll_main_compute57_in[69:6], zll_main_compute57_in[5:3], zll_main_compute57_in[2:0], 3'h5};
  ZLL_Main_compute259  instR7 (zll_main_compute259_inR5[136:73], zll_main_compute259_inR5[72:9], zll_main_compute259_inR5[8:6], zll_main_compute259_inR5[5:3], zll_main_compute259_inR5[2:0], zll_main_compute259_outR5);
  assign zll_main_compute259_inR6 = {zll_main_compute57_in[133:70], zll_main_compute57_in[69:6], zll_main_compute57_in[5:3], zll_main_compute57_in[2:0], 3'h6};
  ZLL_Main_compute259  instR8 (zll_main_compute259_inR6[136:73], zll_main_compute259_inR6[72:9], zll_main_compute259_inR6[8:6], zll_main_compute259_inR6[5:3], zll_main_compute259_inR6[2:0], zll_main_compute259_outR6);
  assign zll_main_compute259_inR7 = {zll_main_compute57_in[133:70], zll_main_compute57_in[69:6], zll_main_compute57_in[5:3], zll_main_compute57_in[2:0], 3'h7};
  ZLL_Main_compute259  instR9 (zll_main_compute259_inR7[136:73], zll_main_compute259_inR7[72:9], zll_main_compute259_inR7[8:6], zll_main_compute259_inR7[5:3], zll_main_compute259_inR7[2:0], zll_main_compute259_outR7);
  assign zll_main_compute124_in = {zll_main_compute191_in[127:64], zll_main_compute191_in[63:0]};
  assign zll_main_compute190_in = {zll_main_compute124_in[127:64], zll_main_compute124_in[63:0]};
  assign zll_main_compute375_in = zll_main_compute190_in[127:0];
  assign zll_main_compute31_in = {zll_main_compute375_in[63:0], zll_main_compute375_in[127:64]};
  assign zll_main_compute148_in = {zll_main_compute31_in[127:64], zll_main_compute31_in[63:0], 3'h1};
  assign zll_main_compute353_in = {zll_main_compute148_in[130:67], zll_main_compute148_in[66:3], zll_main_compute148_in[2:0], 3'h2};
  assign zll_main_compute428_inR1 = {3'h7, zll_main_compute353_in[2:0]};
  ZLL_Main_compute428  instR10 (zll_main_compute428_inR1[5:3], zll_main_compute428_inR1[2:0], zll_main_compute428_outR1);
  assign zll_main_compute70_in = {zll_main_compute353_in[133:70], zll_main_compute353_in[69:6], zll_main_compute353_in[5:3], zll_main_compute353_in[2:0], zll_main_compute428_outR1};
  assign zll_main_compute383_in = {zll_main_compute70_in[2:0], zll_main_compute70_in[72:9], zll_main_compute70_in[8:6], 1'h0};
  ZLL_Main_compute383  instR11 (zll_main_compute383_in[70:68], zll_main_compute383_in[67:4], zll_main_compute383_in[3:1], zll_main_compute383_in[0], zll_main_compute383_out);
  assign zll_main_compute275_in = {zll_main_compute70_in[136:73], zll_main_compute70_in[72:9], zll_main_compute70_in[8:6], zll_main_compute70_in[5:3], zll_main_compute383_out};
  assign zll_main_compute119_in = {zll_main_compute275_in[2:0], zll_main_compute275_in[136:73], zll_main_compute275_in[72:9], zll_main_compute275_in[8:6], zll_main_compute275_in[5:3], 3'h0};
  ZLL_Main_compute119  instR12 (zll_main_compute119_in[139:137], zll_main_compute119_in[136:73], zll_main_compute119_in[72:9], zll_main_compute119_in[8:6], zll_main_compute119_in[5:3], zll_main_compute119_in[2:0], zll_main_compute119_out);
  assign zll_main_compute119_inR1 = {zll_main_compute275_in[2:0], zll_main_compute275_in[136:73], zll_main_compute275_in[72:9], zll_main_compute275_in[8:6], zll_main_compute275_in[5:3], 3'h1};
  ZLL_Main_compute119  instR13 (zll_main_compute119_inR1[139:137], zll_main_compute119_inR1[136:73], zll_main_compute119_inR1[72:9], zll_main_compute119_inR1[8:6], zll_main_compute119_inR1[5:3], zll_main_compute119_inR1[2:0], zll_main_compute119_outR1);
  assign zll_main_compute119_inR2 = {zll_main_compute275_in[2:0], zll_main_compute275_in[136:73], zll_main_compute275_in[72:9], zll_main_compute275_in[8:6], zll_main_compute275_in[5:3], 3'h2};
  ZLL_Main_compute119  instR14 (zll_main_compute119_inR2[139:137], zll_main_compute119_inR2[136:73], zll_main_compute119_inR2[72:9], zll_main_compute119_inR2[8:6], zll_main_compute119_inR2[5:3], zll_main_compute119_inR2[2:0], zll_main_compute119_outR2);
  assign zll_main_compute119_inR3 = {zll_main_compute275_in[2:0], zll_main_compute275_in[136:73], zll_main_compute275_in[72:9], zll_main_compute275_in[8:6], zll_main_compute275_in[5:3], 3'h3};
  ZLL_Main_compute119  instR15 (zll_main_compute119_inR3[139:137], zll_main_compute119_inR3[136:73], zll_main_compute119_inR3[72:9], zll_main_compute119_inR3[8:6], zll_main_compute119_inR3[5:3], zll_main_compute119_inR3[2:0], zll_main_compute119_outR3);
  assign zll_main_compute119_inR4 = {zll_main_compute275_in[2:0], zll_main_compute275_in[136:73], zll_main_compute275_in[72:9], zll_main_compute275_in[8:6], zll_main_compute275_in[5:3], 3'h4};
  ZLL_Main_compute119  instR16 (zll_main_compute119_inR4[139:137], zll_main_compute119_inR4[136:73], zll_main_compute119_inR4[72:9], zll_main_compute119_inR4[8:6], zll_main_compute119_inR4[5:3], zll_main_compute119_inR4[2:0], zll_main_compute119_outR4);
  assign zll_main_compute119_inR5 = {zll_main_compute275_in[2:0], zll_main_compute275_in[136:73], zll_main_compute275_in[72:9], zll_main_compute275_in[8:6], zll_main_compute275_in[5:3], 3'h5};
  ZLL_Main_compute119  instR17 (zll_main_compute119_inR5[139:137], zll_main_compute119_inR5[136:73], zll_main_compute119_inR5[72:9], zll_main_compute119_inR5[8:6], zll_main_compute119_inR5[5:3], zll_main_compute119_inR5[2:0], zll_main_compute119_outR5);
  assign zll_main_compute119_inR6 = {zll_main_compute275_in[2:0], zll_main_compute275_in[136:73], zll_main_compute275_in[72:9], zll_main_compute275_in[8:6], zll_main_compute275_in[5:3], 3'h6};
  ZLL_Main_compute119  instR18 (zll_main_compute119_inR6[139:137], zll_main_compute119_inR6[136:73], zll_main_compute119_inR6[72:9], zll_main_compute119_inR6[8:6], zll_main_compute119_inR6[5:3], zll_main_compute119_inR6[2:0], zll_main_compute119_outR6);
  assign zll_main_compute119_inR7 = {zll_main_compute275_in[2:0], zll_main_compute275_in[136:73], zll_main_compute275_in[72:9], zll_main_compute275_in[8:6], zll_main_compute275_in[5:3], 3'h7};
  ZLL_Main_compute119  instR19 (zll_main_compute119_inR7[139:137], zll_main_compute119_inR7[136:73], zll_main_compute119_inR7[72:9], zll_main_compute119_inR7[8:6], zll_main_compute119_inR7[5:3], zll_main_compute119_inR7[2:0], zll_main_compute119_outR7);
  assign zll_main_compute329_in = {{zll_main_compute259_out, zll_main_compute259_outR1, zll_main_compute259_outR2, zll_main_compute259_outR3, zll_main_compute259_outR4, zll_main_compute259_outR5, zll_main_compute259_outR6, zll_main_compute259_outR7}, {zll_main_compute119_out, zll_main_compute119_outR1, zll_main_compute119_outR2, zll_main_compute119_outR3, zll_main_compute119_outR4, zll_main_compute119_outR5, zll_main_compute119_outR6, zll_main_compute119_outR7}};
  assign zll_main_compute232_in = zll_main_compute329_in[127:0];
  assign zll_main_compute365_in = {zll_main_compute232_in[63:0], zll_main_compute232_in[127:64]};
  assign zll_main_compute254_in = {zll_main_compute365_in[127:64], zll_main_compute365_in[63:0]};
  assign zll_main_compute80_in = zll_main_compute254_in[127:0];
  assign zll_main_compute183_in = {zll_main_compute80_in[127:64], zll_main_compute80_in[63:0], 3'h1};
  assign zll_main_compute422_in = {zll_main_compute183_in[2:0], zll_main_compute183_in[130:67], zll_main_compute183_in[66:3]};
  assign zll_main_compute417_in = {zll_main_compute422_in[130:128], zll_main_compute422_in[127:64], zll_main_compute422_in[63:0], 3'h2};
  assign zll_main_compute428_inR2 = {3'h7, zll_main_compute417_in[2:0]};
  ZLL_Main_compute428  instR20 (zll_main_compute428_inR2[5:3], zll_main_compute428_inR2[2:0], zll_main_compute428_outR2);
  assign zll_main_compute348_in = {zll_main_compute417_in[133:131], zll_main_compute417_in[130:67], zll_main_compute417_in[2:0], zll_main_compute417_in[66:3], zll_main_compute428_outR2};
  assign zll_main_compute6_in = {zll_main_compute348_in[136:134], zll_main_compute348_in[2:0], zll_main_compute348_in[133:70], 1'h0};
  assign zll_main_compute354_inR1 = {zll_main_compute6_in[70:68], zll_main_compute6_in[67:65], 1'h0};
  ZLL_Main_compute354  instR21 (zll_main_compute354_inR1[6:4], zll_main_compute354_inR1[3:1], zll_main_compute354_inR1[0], zll_main_compute354_outR1);
  assign id_inR1 = {zll_main_compute6_in[67:65], zll_main_compute6_in[0]};
  assign zll_main_compute118_in = {zll_main_compute348_in[133:70], zll_main_compute348_in[69:67], zll_main_compute348_in[66:3], (id_inR1[0] == 1'h1) ? id_inR1[3:1] : zll_main_compute354_outR1};
  assign zll_main_compute221_in = {zll_main_compute118_in[2:0], zll_main_compute118_in[133:70], zll_main_compute118_in[69:67], zll_main_compute118_in[66:3], 3'h0};
  ZLL_Main_compute221  instR22 (zll_main_compute221_in[136:134], zll_main_compute221_in[133:70], zll_main_compute221_in[69:67], zll_main_compute221_in[66:3], zll_main_compute221_in[2:0], zll_main_compute221_out);
  assign zll_main_compute221_inR1 = {zll_main_compute118_in[2:0], zll_main_compute118_in[133:70], zll_main_compute118_in[69:67], zll_main_compute118_in[66:3], 3'h1};
  ZLL_Main_compute221  instR23 (zll_main_compute221_inR1[136:134], zll_main_compute221_inR1[133:70], zll_main_compute221_inR1[69:67], zll_main_compute221_inR1[66:3], zll_main_compute221_inR1[2:0], zll_main_compute221_outR1);
  assign zll_main_compute221_inR2 = {zll_main_compute118_in[2:0], zll_main_compute118_in[133:70], zll_main_compute118_in[69:67], zll_main_compute118_in[66:3], 3'h2};
  ZLL_Main_compute221  instR24 (zll_main_compute221_inR2[136:134], zll_main_compute221_inR2[133:70], zll_main_compute221_inR2[69:67], zll_main_compute221_inR2[66:3], zll_main_compute221_inR2[2:0], zll_main_compute221_outR2);
  assign zll_main_compute221_inR3 = {zll_main_compute118_in[2:0], zll_main_compute118_in[133:70], zll_main_compute118_in[69:67], zll_main_compute118_in[66:3], 3'h3};
  ZLL_Main_compute221  instR25 (zll_main_compute221_inR3[136:134], zll_main_compute221_inR3[133:70], zll_main_compute221_inR3[69:67], zll_main_compute221_inR3[66:3], zll_main_compute221_inR3[2:0], zll_main_compute221_outR3);
  assign zll_main_compute221_inR4 = {zll_main_compute118_in[2:0], zll_main_compute118_in[133:70], zll_main_compute118_in[69:67], zll_main_compute118_in[66:3], 3'h4};
  ZLL_Main_compute221  instR26 (zll_main_compute221_inR4[136:134], zll_main_compute221_inR4[133:70], zll_main_compute221_inR4[69:67], zll_main_compute221_inR4[66:3], zll_main_compute221_inR4[2:0], zll_main_compute221_outR4);
  assign zll_main_compute221_inR5 = {zll_main_compute118_in[2:0], zll_main_compute118_in[133:70], zll_main_compute118_in[69:67], zll_main_compute118_in[66:3], 3'h5};
  ZLL_Main_compute221  instR27 (zll_main_compute221_inR5[136:134], zll_main_compute221_inR5[133:70], zll_main_compute221_inR5[69:67], zll_main_compute221_inR5[66:3], zll_main_compute221_inR5[2:0], zll_main_compute221_outR5);
  assign zll_main_compute221_inR6 = {zll_main_compute118_in[2:0], zll_main_compute118_in[133:70], zll_main_compute118_in[69:67], zll_main_compute118_in[66:3], 3'h6};
  ZLL_Main_compute221  instR28 (zll_main_compute221_inR6[136:134], zll_main_compute221_inR6[133:70], zll_main_compute221_inR6[69:67], zll_main_compute221_inR6[66:3], zll_main_compute221_inR6[2:0], zll_main_compute221_outR6);
  assign zll_main_compute221_inR7 = {zll_main_compute118_in[2:0], zll_main_compute118_in[133:70], zll_main_compute118_in[69:67], zll_main_compute118_in[66:3], 3'h7};
  ZLL_Main_compute221  instR29 (zll_main_compute221_inR7[136:134], zll_main_compute221_inR7[133:70], zll_main_compute221_inR7[69:67], zll_main_compute221_inR7[66:3], zll_main_compute221_inR7[2:0], zll_main_compute221_outR7);
  assign zll_main_compute180_in = {zll_main_compute232_in[63:0], zll_main_compute232_in[127:64]};
  assign zll_main_compute20_in = {zll_main_compute180_in[127:64], zll_main_compute180_in[63:0]};
  assign zll_main_compute441_in = zll_main_compute20_in[127:0];
  assign zll_main_compute437_in = {zll_main_compute441_in[63:0], zll_main_compute441_in[127:64]};
  assign zll_main_compute324_in = {zll_main_compute437_in[127:64], zll_main_compute437_in[63:0], 3'h1};
  assign zll_main_compute396_in = {zll_main_compute324_in[130:67], zll_main_compute324_in[2:0], zll_main_compute324_in[66:3]};
  assign zll_main_compute398_in = {zll_main_compute396_in[130:67], zll_main_compute396_in[66:64], zll_main_compute396_in[63:0], 3'h2};
  assign zll_main_compute428_inR3 = {3'h7, zll_main_compute398_in[2:0]};
  ZLL_Main_compute428  instR30 (zll_main_compute428_inR3[5:3], zll_main_compute428_inR3[2:0], zll_main_compute428_outR3);
  assign zll_main_compute407_in = {zll_main_compute398_in[133:70], zll_main_compute398_in[69:67], zll_main_compute398_in[2:0], zll_main_compute398_in[66:3], zll_main_compute428_outR3};
  assign zll_main_compute351_in = {zll_main_compute407_in[2:0], zll_main_compute407_in[72:70], zll_main_compute407_in[66:3], 1'h0};
  assign zll_main_compute321_in = {zll_main_compute351_in[70:68], zll_main_compute351_in[67:65], 1'h0};
  ZLL_Main_compute321  instR31 (zll_main_compute321_in[6:4], zll_main_compute321_in[3:1], zll_main_compute321_in[0], zll_main_compute321_out);
  assign id_inR2 = {zll_main_compute351_in[70:68], zll_main_compute351_in[0]};
  assign zll_main_compute16_in = {zll_main_compute407_in[136:73], zll_main_compute407_in[72:70], zll_main_compute407_in[69:67], zll_main_compute407_in[66:3], (id_inR2[0] == 1'h1) ? id_inR2[3:1] : zll_main_compute321_out};
  assign zll_main_compute28_in = {zll_main_compute16_in[136:73], zll_main_compute16_in[72:70], zll_main_compute16_in[69:67], zll_main_compute16_in[2:0], zll_main_compute16_in[66:3], 3'h0};
  ZLL_Main_compute28  instR32 (zll_main_compute28_in[139:76], zll_main_compute28_in[75:73], zll_main_compute28_in[72:70], zll_main_compute28_in[69:67], zll_main_compute28_in[66:3], zll_main_compute28_in[2:0], zll_main_compute28_out);
  assign zll_main_compute28_inR1 = {zll_main_compute16_in[136:73], zll_main_compute16_in[72:70], zll_main_compute16_in[69:67], zll_main_compute16_in[2:0], zll_main_compute16_in[66:3], 3'h1};
  ZLL_Main_compute28  instR33 (zll_main_compute28_inR1[139:76], zll_main_compute28_inR1[75:73], zll_main_compute28_inR1[72:70], zll_main_compute28_inR1[69:67], zll_main_compute28_inR1[66:3], zll_main_compute28_inR1[2:0], zll_main_compute28_outR1);
  assign zll_main_compute28_inR2 = {zll_main_compute16_in[136:73], zll_main_compute16_in[72:70], zll_main_compute16_in[69:67], zll_main_compute16_in[2:0], zll_main_compute16_in[66:3], 3'h2};
  ZLL_Main_compute28  instR34 (zll_main_compute28_inR2[139:76], zll_main_compute28_inR2[75:73], zll_main_compute28_inR2[72:70], zll_main_compute28_inR2[69:67], zll_main_compute28_inR2[66:3], zll_main_compute28_inR2[2:0], zll_main_compute28_outR2);
  assign zll_main_compute28_inR3 = {zll_main_compute16_in[136:73], zll_main_compute16_in[72:70], zll_main_compute16_in[69:67], zll_main_compute16_in[2:0], zll_main_compute16_in[66:3], 3'h3};
  ZLL_Main_compute28  instR35 (zll_main_compute28_inR3[139:76], zll_main_compute28_inR3[75:73], zll_main_compute28_inR3[72:70], zll_main_compute28_inR3[69:67], zll_main_compute28_inR3[66:3], zll_main_compute28_inR3[2:0], zll_main_compute28_outR3);
  assign zll_main_compute28_inR4 = {zll_main_compute16_in[136:73], zll_main_compute16_in[72:70], zll_main_compute16_in[69:67], zll_main_compute16_in[2:0], zll_main_compute16_in[66:3], 3'h4};
  ZLL_Main_compute28  instR36 (zll_main_compute28_inR4[139:76], zll_main_compute28_inR4[75:73], zll_main_compute28_inR4[72:70], zll_main_compute28_inR4[69:67], zll_main_compute28_inR4[66:3], zll_main_compute28_inR4[2:0], zll_main_compute28_outR4);
  assign zll_main_compute28_inR5 = {zll_main_compute16_in[136:73], zll_main_compute16_in[72:70], zll_main_compute16_in[69:67], zll_main_compute16_in[2:0], zll_main_compute16_in[66:3], 3'h5};
  ZLL_Main_compute28  instR37 (zll_main_compute28_inR5[139:76], zll_main_compute28_inR5[75:73], zll_main_compute28_inR5[72:70], zll_main_compute28_inR5[69:67], zll_main_compute28_inR5[66:3], zll_main_compute28_inR5[2:0], zll_main_compute28_outR5);
  assign zll_main_compute28_inR6 = {zll_main_compute16_in[136:73], zll_main_compute16_in[72:70], zll_main_compute16_in[69:67], zll_main_compute16_in[2:0], zll_main_compute16_in[66:3], 3'h6};
  ZLL_Main_compute28  instR38 (zll_main_compute28_inR6[139:76], zll_main_compute28_inR6[75:73], zll_main_compute28_inR6[72:70], zll_main_compute28_inR6[69:67], zll_main_compute28_inR6[66:3], zll_main_compute28_inR6[2:0], zll_main_compute28_outR6);
  assign zll_main_compute28_inR7 = {zll_main_compute16_in[136:73], zll_main_compute16_in[72:70], zll_main_compute16_in[69:67], zll_main_compute16_in[2:0], zll_main_compute16_in[66:3], 3'h7};
  ZLL_Main_compute28  instR39 (zll_main_compute28_inR7[139:76], zll_main_compute28_inR7[75:73], zll_main_compute28_inR7[72:70], zll_main_compute28_inR7[69:67], zll_main_compute28_inR7[66:3], zll_main_compute28_inR7[2:0], zll_main_compute28_outR7);
  assign zll_main_compute97_in = {{zll_main_compute221_out, zll_main_compute221_outR1, zll_main_compute221_outR2, zll_main_compute221_outR3, zll_main_compute221_outR4, zll_main_compute221_outR5, zll_main_compute221_outR6, zll_main_compute221_outR7}, {zll_main_compute28_out, zll_main_compute28_outR1, zll_main_compute28_outR2, zll_main_compute28_outR3, zll_main_compute28_outR4, zll_main_compute28_outR5, zll_main_compute28_outR6, zll_main_compute28_outR7}};
  assign zll_main_compute357_in = zll_main_compute97_in[127:0];
  assign zll_main_compute293_in = {zll_main_compute357_in[127:64], zll_main_compute357_in[63:0]};
  assign zll_main_compute371_in = {zll_main_compute293_in[127:64], zll_main_compute293_in[63:0]};
  assign zll_main_compute160_in = zll_main_compute371_in[127:0];
  assign zll_main_compute279_in = {zll_main_compute160_in[63:0], zll_main_compute160_in[127:64]};
  assign zll_main_compute178_in = {zll_main_compute279_in[127:64], zll_main_compute279_in[63:0], 3'h1};
  assign zll_main_compute261_in = {zll_main_compute178_in[130:67], zll_main_compute178_in[66:3], zll_main_compute178_in[2:0], 3'h2};
  assign zll_main_compute198_in = {zll_main_compute261_in[133:70], zll_main_compute261_in[2:0], zll_main_compute261_in[69:6], zll_main_compute261_in[5:3], 3'h0};
  ZLL_Main_compute198  instR40 (zll_main_compute198_in[136:73], zll_main_compute198_in[72:70], zll_main_compute198_in[69:6], zll_main_compute198_in[5:3], zll_main_compute198_in[2:0], zll_main_compute198_out);
  assign zll_main_compute198_inR1 = {zll_main_compute261_in[133:70], zll_main_compute261_in[2:0], zll_main_compute261_in[69:6], zll_main_compute261_in[5:3], 3'h1};
  ZLL_Main_compute198  instR41 (zll_main_compute198_inR1[136:73], zll_main_compute198_inR1[72:70], zll_main_compute198_inR1[69:6], zll_main_compute198_inR1[5:3], zll_main_compute198_inR1[2:0], zll_main_compute198_outR1);
  assign zll_main_compute198_inR2 = {zll_main_compute261_in[133:70], zll_main_compute261_in[2:0], zll_main_compute261_in[69:6], zll_main_compute261_in[5:3], 3'h2};
  ZLL_Main_compute198  instR42 (zll_main_compute198_inR2[136:73], zll_main_compute198_inR2[72:70], zll_main_compute198_inR2[69:6], zll_main_compute198_inR2[5:3], zll_main_compute198_inR2[2:0], zll_main_compute198_outR2);
  assign zll_main_compute198_inR3 = {zll_main_compute261_in[133:70], zll_main_compute261_in[2:0], zll_main_compute261_in[69:6], zll_main_compute261_in[5:3], 3'h3};
  ZLL_Main_compute198  instR43 (zll_main_compute198_inR3[136:73], zll_main_compute198_inR3[72:70], zll_main_compute198_inR3[69:6], zll_main_compute198_inR3[5:3], zll_main_compute198_inR3[2:0], zll_main_compute198_outR3);
  assign zll_main_compute198_inR4 = {zll_main_compute261_in[133:70], zll_main_compute261_in[2:0], zll_main_compute261_in[69:6], zll_main_compute261_in[5:3], 3'h4};
  ZLL_Main_compute198  instR44 (zll_main_compute198_inR4[136:73], zll_main_compute198_inR4[72:70], zll_main_compute198_inR4[69:6], zll_main_compute198_inR4[5:3], zll_main_compute198_inR4[2:0], zll_main_compute198_outR4);
  assign zll_main_compute198_inR5 = {zll_main_compute261_in[133:70], zll_main_compute261_in[2:0], zll_main_compute261_in[69:6], zll_main_compute261_in[5:3], 3'h5};
  ZLL_Main_compute198  instR45 (zll_main_compute198_inR5[136:73], zll_main_compute198_inR5[72:70], zll_main_compute198_inR5[69:6], zll_main_compute198_inR5[5:3], zll_main_compute198_inR5[2:0], zll_main_compute198_outR5);
  assign zll_main_compute198_inR6 = {zll_main_compute261_in[133:70], zll_main_compute261_in[2:0], zll_main_compute261_in[69:6], zll_main_compute261_in[5:3], 3'h6};
  ZLL_Main_compute198  instR46 (zll_main_compute198_inR6[136:73], zll_main_compute198_inR6[72:70], zll_main_compute198_inR6[69:6], zll_main_compute198_inR6[5:3], zll_main_compute198_inR6[2:0], zll_main_compute198_outR6);
  assign zll_main_compute198_inR7 = {zll_main_compute261_in[133:70], zll_main_compute261_in[2:0], zll_main_compute261_in[69:6], zll_main_compute261_in[5:3], 3'h7};
  ZLL_Main_compute198  instR47 (zll_main_compute198_inR7[136:73], zll_main_compute198_inR7[72:70], zll_main_compute198_inR7[69:6], zll_main_compute198_inR7[5:3], zll_main_compute198_inR7[2:0], zll_main_compute198_outR7);
  assign zll_main_compute286_in = {zll_main_compute357_in[127:64], zll_main_compute357_in[63:0]};
  assign zll_main_compute127_in = {zll_main_compute286_in[127:64], zll_main_compute286_in[63:0]};
  assign zll_main_compute399_in = zll_main_compute127_in[127:0];
  assign zll_main_compute243_in = {zll_main_compute399_in[127:64], zll_main_compute399_in[63:0], 3'h1};
  assign zll_main_compute55_in = {zll_main_compute243_in[130:67], zll_main_compute243_in[66:3], zll_main_compute243_in[2:0], 3'h2};
  assign zll_main_compute428_inR4 = {3'h7, zll_main_compute55_in[2:0]};
  ZLL_Main_compute428  instR48 (zll_main_compute428_inR4[5:3], zll_main_compute428_inR4[2:0], zll_main_compute428_outR4);
  assign zll_main_compute96_in = {zll_main_compute55_in[2:0], zll_main_compute55_in[133:70], zll_main_compute55_in[69:6], zll_main_compute55_in[5:3], zll_main_compute428_outR4};
  assign zll_main_compute383_inR1 = {zll_main_compute96_in[2:0], zll_main_compute96_in[133:70], zll_main_compute96_in[5:3], 1'h0};
  ZLL_Main_compute383  instR49 (zll_main_compute383_inR1[70:68], zll_main_compute383_inR1[67:4], zll_main_compute383_inR1[3:1], zll_main_compute383_inR1[0], zll_main_compute383_outR1);
  assign zll_main_compute406_in = {zll_main_compute96_in[136:134], zll_main_compute96_in[133:70], zll_main_compute96_in[69:6], zll_main_compute96_in[5:3], zll_main_compute383_outR1};
  assign zll_main_compute141_in = {zll_main_compute406_in[136:134], zll_main_compute406_in[2:0], zll_main_compute406_in[133:70], zll_main_compute406_in[69:6], zll_main_compute406_in[5:3], 3'h0};
  ZLL_Main_compute141  instR50 (zll_main_compute141_in[139:137], zll_main_compute141_in[136:134], zll_main_compute141_in[133:70], zll_main_compute141_in[69:6], zll_main_compute141_in[5:3], zll_main_compute141_in[2:0], zll_main_compute141_out);
  assign zll_main_compute141_inR1 = {zll_main_compute406_in[136:134], zll_main_compute406_in[2:0], zll_main_compute406_in[133:70], zll_main_compute406_in[69:6], zll_main_compute406_in[5:3], 3'h1};
  ZLL_Main_compute141  instR51 (zll_main_compute141_inR1[139:137], zll_main_compute141_inR1[136:134], zll_main_compute141_inR1[133:70], zll_main_compute141_inR1[69:6], zll_main_compute141_inR1[5:3], zll_main_compute141_inR1[2:0], zll_main_compute141_outR1);
  assign zll_main_compute141_inR2 = {zll_main_compute406_in[136:134], zll_main_compute406_in[2:0], zll_main_compute406_in[133:70], zll_main_compute406_in[69:6], zll_main_compute406_in[5:3], 3'h2};
  ZLL_Main_compute141  instR52 (zll_main_compute141_inR2[139:137], zll_main_compute141_inR2[136:134], zll_main_compute141_inR2[133:70], zll_main_compute141_inR2[69:6], zll_main_compute141_inR2[5:3], zll_main_compute141_inR2[2:0], zll_main_compute141_outR2);
  assign zll_main_compute141_inR3 = {zll_main_compute406_in[136:134], zll_main_compute406_in[2:0], zll_main_compute406_in[133:70], zll_main_compute406_in[69:6], zll_main_compute406_in[5:3], 3'h3};
  ZLL_Main_compute141  instR53 (zll_main_compute141_inR3[139:137], zll_main_compute141_inR3[136:134], zll_main_compute141_inR3[133:70], zll_main_compute141_inR3[69:6], zll_main_compute141_inR3[5:3], zll_main_compute141_inR3[2:0], zll_main_compute141_outR3);
  assign zll_main_compute141_inR4 = {zll_main_compute406_in[136:134], zll_main_compute406_in[2:0], zll_main_compute406_in[133:70], zll_main_compute406_in[69:6], zll_main_compute406_in[5:3], 3'h4};
  ZLL_Main_compute141  instR54 (zll_main_compute141_inR4[139:137], zll_main_compute141_inR4[136:134], zll_main_compute141_inR4[133:70], zll_main_compute141_inR4[69:6], zll_main_compute141_inR4[5:3], zll_main_compute141_inR4[2:0], zll_main_compute141_outR4);
  assign zll_main_compute141_inR5 = {zll_main_compute406_in[136:134], zll_main_compute406_in[2:0], zll_main_compute406_in[133:70], zll_main_compute406_in[69:6], zll_main_compute406_in[5:3], 3'h5};
  ZLL_Main_compute141  instR55 (zll_main_compute141_inR5[139:137], zll_main_compute141_inR5[136:134], zll_main_compute141_inR5[133:70], zll_main_compute141_inR5[69:6], zll_main_compute141_inR5[5:3], zll_main_compute141_inR5[2:0], zll_main_compute141_outR5);
  assign zll_main_compute141_inR6 = {zll_main_compute406_in[136:134], zll_main_compute406_in[2:0], zll_main_compute406_in[133:70], zll_main_compute406_in[69:6], zll_main_compute406_in[5:3], 3'h6};
  ZLL_Main_compute141  instR56 (zll_main_compute141_inR6[139:137], zll_main_compute141_inR6[136:134], zll_main_compute141_inR6[133:70], zll_main_compute141_inR6[69:6], zll_main_compute141_inR6[5:3], zll_main_compute141_inR6[2:0], zll_main_compute141_outR6);
  assign zll_main_compute141_inR7 = {zll_main_compute406_in[136:134], zll_main_compute406_in[2:0], zll_main_compute406_in[133:70], zll_main_compute406_in[69:6], zll_main_compute406_in[5:3], 3'h7};
  ZLL_Main_compute141  instR57 (zll_main_compute141_inR7[139:137], zll_main_compute141_inR7[136:134], zll_main_compute141_inR7[133:70], zll_main_compute141_inR7[69:6], zll_main_compute141_inR7[5:3], zll_main_compute141_inR7[2:0], zll_main_compute141_outR7);
  assign zll_main_compute442_in = {{zll_main_compute198_out, zll_main_compute198_outR1, zll_main_compute198_outR2, zll_main_compute198_outR3, zll_main_compute198_outR4, zll_main_compute198_outR5, zll_main_compute198_outR6, zll_main_compute198_outR7}, {zll_main_compute141_out, zll_main_compute141_outR1, zll_main_compute141_outR2, zll_main_compute141_outR3, zll_main_compute141_outR4, zll_main_compute141_outR5, zll_main_compute141_outR6, zll_main_compute141_outR7}};
  assign id_inR3 = zll_main_compute442_in[127:0];
  assign zll_main_loop1_in = {1'h0, {id_inR3[127:64], id_inR3[63:0]}};
  assign zll_main_loop2_in = zll_main_loop1_in[128:0];
  assign {__continue, __out0, __out1} = {1'h1, zll_main_loop2_in[127:0]};
endmodule

module ZLL_Main_compute450 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  output logic [2:0] res);
  logic [5:0] zll_main_compute328_in;
  logic [5:0] zll_main_compute423_in;
  logic [2:0] resize_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR2;
  assign zll_main_compute328_in = {arg0, arg1};
  assign zll_main_compute423_in = zll_main_compute328_in[5:0];
  assign resize_in = zll_main_compute423_in[5:3];
  assign resize_inR1 = zll_main_compute423_in[2:0];
  assign binop_in = {128'(resize_in[2:0]), 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] + binop_in[127:0], 128'h8};
  assign resize_inR2 = binop_inR1[255:128] % binop_inR1[127:0];
  assign res = resize_inR2[2:0];
endmodule

module ZLL_Main_compute447 (input logic [2:0] arg0,
  output logic [0:0] res);
  logic [2:0] resize_in;
  logic [127:0] zll_main_compute368_in;
  logic [127:0] resize_inR1;
  logic [0:0] msbit_in;
  logic [0:0] rewire_prelude_not_in;
  logic [1:0] zll_rewire_prelude_not2_in;
  logic [0:0] lit_in;
  assign resize_in = arg0;
  assign zll_main_compute368_in = 128'(resize_in[2:0]);
  assign resize_inR1 = zll_main_compute368_in[127:0];
  assign msbit_in = resize_inR1[0];
  assign rewire_prelude_not_in = msbit_in[0];
  assign zll_rewire_prelude_not2_in = {rewire_prelude_not_in[0], rewire_prelude_not_in[0]};
  assign lit_in = zll_rewire_prelude_not2_in[0];
  assign res = (lit_in[0] == 1'h1) ? 1'h0 : 1'h1;
endmodule

module ZLL_Main_compute428 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  output logic [2:0] res);
  logic [5:0] zll_main_compute436_in;
  logic [5:0] zll_main_compute408_in;
  logic [2:0] resize_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR2;
  assign zll_main_compute436_in = {arg0, arg1};
  assign zll_main_compute408_in = zll_main_compute436_in[5:0];
  assign resize_in = zll_main_compute408_in[5:3];
  assign resize_inR1 = zll_main_compute408_in[2:0];
  assign binop_in = {128'(resize_in[2:0]), 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] / binop_in[127:0], 128'h8};
  assign resize_inR2 = binop_inR1[255:128] % binop_inR1[127:0];
  assign res = resize_inR2[2:0];
endmodule

module ZLL_Main_compute412 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  output logic [0:0] res);
  logic [5:0] zll_main_compute393_in;
  logic [5:0] zll_main_compute444_in;
  logic [2:0] resize_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  assign zll_main_compute393_in = {arg0, arg1};
  assign zll_main_compute444_in = zll_main_compute393_in[5:0];
  assign resize_in = zll_main_compute444_in[5:3];
  assign resize_inR1 = zll_main_compute444_in[2:0];
  assign binop_in = {128'(resize_in[2:0]), 128'(resize_inR1[2:0])};
  assign res = binop_in[255:128] < binop_in[127:0];
endmodule

module ZLL_Main_compute383 (input logic [2:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  input logic [0:0] arg3,
  output logic [2:0] res);
  logic [6:0] zll_main_compute321_in;
  logic [2:0] zll_main_compute321_out;
  logic [3:0] id_in;
  assign zll_main_compute321_in = {arg0, arg2, 1'h0};
  ZLL_Main_compute321  inst (zll_main_compute321_in[6:4], zll_main_compute321_in[3:1], zll_main_compute321_in[0], zll_main_compute321_out);
  assign id_in = {arg0, arg3};
  assign res = (id_in[0] == 1'h1) ? id_in[3:1] : zll_main_compute321_out;
endmodule

module ZLL_Main_compute373 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  output logic [2:0] res);
  logic [5:0] zll_main_compute448_in;
  logic [5:0] zll_main_compute378_in;
  logic [2:0] resize_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR2;
  assign zll_main_compute448_in = {arg0, arg1};
  assign zll_main_compute378_in = zll_main_compute448_in[5:0];
  assign resize_in = zll_main_compute378_in[5:3];
  assign resize_inR1 = zll_main_compute378_in[2:0];
  assign binop_in = {128'(resize_in[2:0]), 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h8};
  assign resize_inR2 = binop_inR1[255:128] % binop_inR1[127:0];
  assign res = resize_inR2[2:0];
endmodule

module ZLL_Main_compute354 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  input logic [0:0] arg2,
  output logic [2:0] res);
  logic [6:0] zll_main_compute376_in;
  logic [5:0] zll_main_compute450_in;
  logic [2:0] zll_main_compute450_out;
  assign zll_main_compute376_in = {arg0, arg1, arg2};
  assign zll_main_compute450_in = {zll_main_compute376_in[3:1], zll_main_compute376_in[6:4]};
  ZLL_Main_compute450  inst (zll_main_compute450_in[5:3], zll_main_compute450_in[2:0], zll_main_compute450_out);
  assign res = zll_main_compute450_out;
endmodule

module ZLL_Main_compute326 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  output logic [2:0] res);
  logic [5:0] zll_main_compute433_in;
  logic [5:0] zll_main_compute451_in;
  logic [2:0] resize_in;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [127:0] resize_inR2;
  assign zll_main_compute433_in = {arg0, arg1};
  assign zll_main_compute451_in = zll_main_compute433_in[5:0];
  assign resize_in = zll_main_compute451_in[5:3];
  assign resize_inR1 = zll_main_compute451_in[2:0];
  assign binop_in = {128'(resize_in[2:0]), 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] * binop_in[127:0], 128'h8};
  assign resize_inR2 = binop_inR1[255:128] % binop_inR1[127:0];
  assign res = resize_inR2[2:0];
endmodule

module ZLL_Main_compute321 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  input logic [0:0] arg2,
  output logic [2:0] res);
  logic [6:0] zll_main_compute294_in;
  logic [5:0] zll_main_compute450_in;
  logic [2:0] zll_main_compute450_out;
  assign zll_main_compute294_in = {arg0, arg1, arg2};
  assign zll_main_compute450_in = {zll_main_compute294_in[6:4], zll_main_compute294_in[3:1]};
  ZLL_Main_compute450  inst (zll_main_compute450_in[5:3], zll_main_compute450_in[2:0], zll_main_compute450_out);
  assign res = zll_main_compute450_out;
endmodule

module ZLL_Main_compute259 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  input logic [2:0] arg3,
  input logic [2:0] arg4,
  output logic [7:0] res);
  logic [5:0] zll_main_compute412_in;
  logic [0:0] zll_main_compute412_out;
  logic [137:0] zll_main_compute138_in;
  logic [5:0] zll_main_compute412_inR1;
  logic [0:0] zll_main_compute412_outR1;
  logic [73:0] zll_main_compute33_in;
  logic [73:0] zll_main_compute360_in;
  logic [63:0] resize_in;
  logic [5:0] zll_main_compute373_in;
  logic [2:0] zll_main_compute373_out;
  logic [5:0] zll_main_compute326_in;
  logic [2:0] zll_main_compute326_out;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR2;
  logic [70:0] zll_main_compute253_in;
  logic [63:0] resize_inR3;
  logic [5:0] zll_main_compute326_inR1;
  logic [2:0] zll_main_compute326_outR1;
  logic [2:0] resize_inR4;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR5;
  assign zll_main_compute412_in = {arg4, arg3};
  ZLL_Main_compute412  inst (zll_main_compute412_in[5:3], zll_main_compute412_in[2:0], zll_main_compute412_out);
  assign zll_main_compute138_in = {arg0, arg1, arg2, arg4, arg3, zll_main_compute412_out};
  assign zll_main_compute412_inR1 = {zll_main_compute138_in[6:4], zll_main_compute138_in[3:1]};
  ZLL_Main_compute412  instR1 (zll_main_compute412_inR1[5:3], zll_main_compute412_inR1[2:0], zll_main_compute412_outR1);
  assign zll_main_compute33_in = {zll_main_compute138_in[73:10], zll_main_compute138_in[9:7], zll_main_compute138_in[6:4], zll_main_compute138_in[3:1], zll_main_compute412_outR1};
  assign zll_main_compute360_in = {zll_main_compute33_in[73:10], zll_main_compute33_in[9:7], zll_main_compute33_in[6:4], zll_main_compute33_in[3:1], zll_main_compute33_in[0]};
  assign resize_in = zll_main_compute360_in[73:10];
  assign zll_main_compute373_in = {zll_main_compute360_in[6:4], zll_main_compute360_in[3:1]};
  ZLL_Main_compute373  instR2 (zll_main_compute373_in[5:3], zll_main_compute373_in[2:0], zll_main_compute373_out);
  assign zll_main_compute326_in = {zll_main_compute373_out, zll_main_compute360_in[9:7]};
  ZLL_Main_compute326  instR3 (zll_main_compute326_in[5:3], zll_main_compute326_in[2:0], zll_main_compute326_out);
  assign resize_inR1 = zll_main_compute326_out;
  assign binop_in = {128'h8, 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h8};
  assign binop_inR3 = {128'(resize_in[63:0]), binop_inR2[255:128] * binop_inR2[127:0]};
  assign resize_inR2 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign zll_main_compute253_in = {zll_main_compute138_in[137:74], zll_main_compute138_in[9:7], zll_main_compute138_in[6:4], zll_main_compute138_in[0]};
  assign resize_inR3 = zll_main_compute253_in[70:7];
  assign zll_main_compute326_inR1 = {zll_main_compute253_in[3:1], zll_main_compute253_in[6:4]};
  ZLL_Main_compute326  instR4 (zll_main_compute326_inR1[5:3], zll_main_compute326_inR1[2:0], zll_main_compute326_outR1);
  assign resize_inR4 = zll_main_compute326_outR1;
  assign binop_inR4 = {128'h8, 128'(resize_inR4[2:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h8};
  assign binop_inR7 = {128'(resize_inR3[63:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR5 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign res = (zll_main_compute253_in[0] == 1'h1) ? resize_inR5[7:0] : resize_inR2[7:0];
endmodule

module ZLL_Main_compute221 (input logic [2:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  input logic [63:0] arg3,
  input logic [2:0] arg4,
  output logic [7:0] res);
  logic [5:0] zll_main_compute412_in;
  logic [0:0] zll_main_compute412_out;
  logic [137:0] zll_main_compute258_in;
  logic [5:0] zll_main_compute412_inR1;
  logic [0:0] zll_main_compute412_outR1;
  logic [73:0] zll_main_compute155_in;
  logic [73:0] zll_main_compute331_in;
  logic [63:0] resize_in;
  logic [5:0] zll_main_compute373_in;
  logic [2:0] zll_main_compute373_out;
  logic [5:0] zll_main_compute326_in;
  logic [2:0] zll_main_compute326_out;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR2;
  logic [70:0] zll_main_compute318_in;
  logic [63:0] resize_inR3;
  logic [5:0] zll_main_compute326_inR1;
  logic [2:0] zll_main_compute326_outR1;
  logic [2:0] resize_inR4;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR5;
  assign zll_main_compute412_in = {arg4, arg0};
  ZLL_Main_compute412  inst (zll_main_compute412_in[5:3], zll_main_compute412_in[2:0], zll_main_compute412_out);
  assign zll_main_compute258_in = {arg0, arg4, arg1, arg2, arg3, zll_main_compute412_out};
  assign zll_main_compute412_inR1 = {zll_main_compute258_in[134:132], zll_main_compute258_in[137:135]};
  ZLL_Main_compute412  instR1 (zll_main_compute412_inR1[5:3], zll_main_compute412_inR1[2:0], zll_main_compute412_outR1);
  assign zll_main_compute155_in = {zll_main_compute258_in[137:135], zll_main_compute258_in[134:132], zll_main_compute258_in[67:65], zll_main_compute258_in[64:1], zll_main_compute412_outR1};
  assign zll_main_compute331_in = {zll_main_compute155_in[73:71], zll_main_compute155_in[70:68], zll_main_compute155_in[67:65], zll_main_compute155_in[64:1], zll_main_compute155_in[0]};
  assign resize_in = zll_main_compute331_in[64:1];
  assign zll_main_compute373_in = {zll_main_compute331_in[70:68], zll_main_compute331_in[73:71]};
  ZLL_Main_compute373  instR2 (zll_main_compute373_in[5:3], zll_main_compute373_in[2:0], zll_main_compute373_out);
  assign zll_main_compute326_in = {zll_main_compute373_out, zll_main_compute331_in[67:65]};
  ZLL_Main_compute326  instR3 (zll_main_compute326_in[5:3], zll_main_compute326_in[2:0], zll_main_compute326_out);
  assign resize_inR1 = zll_main_compute326_out;
  assign binop_in = {128'h8, 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h8};
  assign binop_inR3 = {128'(resize_in[63:0]), binop_inR2[255:128] * binop_inR2[127:0]};
  assign resize_inR2 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign zll_main_compute318_in = {zll_main_compute258_in[134:132], zll_main_compute258_in[131:68], zll_main_compute258_in[67:65], zll_main_compute258_in[0]};
  assign resize_inR3 = zll_main_compute318_in[67:4];
  assign zll_main_compute326_inR1 = {zll_main_compute318_in[70:68], zll_main_compute318_in[3:1]};
  ZLL_Main_compute326  instR4 (zll_main_compute326_inR1[5:3], zll_main_compute326_inR1[2:0], zll_main_compute326_outR1);
  assign resize_inR4 = zll_main_compute326_outR1;
  assign binop_inR4 = {128'h8, 128'(resize_inR4[2:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h8};
  assign binop_inR7 = {128'(resize_inR3[63:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR5 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign res = (zll_main_compute318_in[0] == 1'h1) ? resize_inR5[7:0] : resize_inR2[7:0];
endmodule

module ZLL_Main_compute198 (input logic [63:0] arg0,
  input logic [2:0] arg1,
  input logic [63:0] arg2,
  input logic [2:0] arg3,
  input logic [2:0] arg4,
  output logic [7:0] res);
  logic [2:0] zll_main_compute447_in;
  logic [0:0] zll_main_compute447_out;
  logic [137:0] zll_main_compute319_in;
  logic [2:0] zll_main_compute447_inR1;
  logic [0:0] zll_main_compute447_outR1;
  logic [73:0] zll_main_compute391_in;
  logic [73:0] zll_main_compute305_in;
  logic [63:0] resize_in;
  logic [5:0] zll_main_compute373_in;
  logic [2:0] zll_main_compute373_out;
  logic [5:0] zll_main_compute428_in;
  logic [2:0] zll_main_compute428_out;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR2;
  logic [70:0] zll_main_compute435_in;
  logic [63:0] resize_inR3;
  logic [5:0] zll_main_compute428_inR1;
  logic [2:0] zll_main_compute428_outR1;
  logic [2:0] resize_inR4;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR5;
  assign zll_main_compute447_in = arg4;
  ZLL_Main_compute447  inst (zll_main_compute447_in[2:0], zll_main_compute447_out);
  assign zll_main_compute319_in = {arg0, arg1, arg2, arg3, arg4, zll_main_compute447_out};
  assign zll_main_compute447_inR1 = zll_main_compute319_in[3:1];
  ZLL_Main_compute447  instR1 (zll_main_compute447_inR1[2:0], zll_main_compute447_outR1);
  assign zll_main_compute391_in = {zll_main_compute319_in[137:74], zll_main_compute319_in[73:71], zll_main_compute319_in[6:4], zll_main_compute319_in[3:1], zll_main_compute447_outR1};
  assign zll_main_compute305_in = {zll_main_compute391_in[73:10], zll_main_compute391_in[9:7], zll_main_compute391_in[6:4], zll_main_compute391_in[3:1], zll_main_compute391_in[0]};
  assign resize_in = zll_main_compute305_in[73:10];
  assign zll_main_compute373_in = {zll_main_compute305_in[3:1], zll_main_compute305_in[6:4]};
  ZLL_Main_compute373  instR2 (zll_main_compute373_in[5:3], zll_main_compute373_in[2:0], zll_main_compute373_out);
  assign zll_main_compute428_in = {zll_main_compute373_out, zll_main_compute305_in[9:7]};
  ZLL_Main_compute428  instR3 (zll_main_compute428_in[5:3], zll_main_compute428_in[2:0], zll_main_compute428_out);
  assign resize_inR1 = zll_main_compute428_out;
  assign binop_in = {128'h8, 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h8};
  assign binop_inR3 = {128'(resize_in[63:0]), binop_inR2[255:128] * binop_inR2[127:0]};
  assign resize_inR2 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign zll_main_compute435_in = {zll_main_compute319_in[73:71], zll_main_compute319_in[70:7], zll_main_compute319_in[3:1], zll_main_compute319_in[0]};
  assign resize_inR3 = zll_main_compute435_in[67:4];
  assign zll_main_compute428_inR1 = {zll_main_compute435_in[3:1], zll_main_compute435_in[70:68]};
  ZLL_Main_compute428  instR4 (zll_main_compute428_inR1[5:3], zll_main_compute428_inR1[2:0], zll_main_compute428_outR1);
  assign resize_inR4 = zll_main_compute428_outR1;
  assign binop_inR4 = {128'h8, 128'(resize_inR4[2:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h8};
  assign binop_inR7 = {128'(resize_inR3[63:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR5 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign res = (zll_main_compute435_in[0] == 1'h1) ? resize_inR5[7:0] : resize_inR2[7:0];
endmodule

module ZLL_Main_compute141 (input logic [2:0] arg0,
  input logic [2:0] arg1,
  input logic [63:0] arg2,
  input logic [63:0] arg3,
  input logic [2:0] arg4,
  input logic [2:0] arg5,
  output logic [7:0] res);
  logic [2:0] zll_main_compute447_in;
  logic [0:0] zll_main_compute447_out;
  logic [140:0] zll_main_compute225_in;
  logic [2:0] zll_main_compute447_inR1;
  logic [0:0] zll_main_compute447_outR1;
  logic [76:0] zll_main_compute157_in;
  logic [76:0] zll_main_compute228_in;
  logic [63:0] resize_in;
  logic [5:0] zll_main_compute373_in;
  logic [2:0] zll_main_compute373_out;
  logic [5:0] zll_main_compute428_in;
  logic [2:0] zll_main_compute428_out;
  logic [5:0] zll_main_compute450_in;
  logic [2:0] zll_main_compute450_out;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR2;
  logic [73:0] zll_main_compute10_in;
  logic [63:0] resize_inR3;
  logic [5:0] zll_main_compute428_inR1;
  logic [2:0] zll_main_compute428_outR1;
  logic [5:0] zll_main_compute450_inR1;
  logic [2:0] zll_main_compute450_outR1;
  logic [2:0] resize_inR4;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR5;
  assign zll_main_compute447_in = arg5;
  ZLL_Main_compute447  inst (zll_main_compute447_in[2:0], zll_main_compute447_out);
  assign zll_main_compute225_in = {arg0, arg1, arg2, arg3, arg4, arg5, zll_main_compute447_out};
  assign zll_main_compute447_inR1 = zll_main_compute225_in[3:1];
  ZLL_Main_compute447  instR1 (zll_main_compute447_inR1[2:0], zll_main_compute447_outR1);
  assign zll_main_compute157_in = {zll_main_compute225_in[140:138], zll_main_compute225_in[137:135], zll_main_compute225_in[70:7], zll_main_compute225_in[6:4], zll_main_compute225_in[3:1], zll_main_compute447_outR1};
  assign zll_main_compute228_in = {zll_main_compute157_in[76:74], zll_main_compute157_in[73:71], zll_main_compute157_in[70:7], zll_main_compute157_in[6:4], zll_main_compute157_in[3:1], zll_main_compute157_in[0]};
  assign resize_in = zll_main_compute228_in[70:7];
  assign zll_main_compute373_in = {zll_main_compute228_in[3:1], zll_main_compute228_in[6:4]};
  ZLL_Main_compute373  instR2 (zll_main_compute373_in[5:3], zll_main_compute373_in[2:0], zll_main_compute373_out);
  assign zll_main_compute428_in = {zll_main_compute373_out, zll_main_compute228_in[76:74]};
  ZLL_Main_compute428  instR3 (zll_main_compute428_in[5:3], zll_main_compute428_in[2:0], zll_main_compute428_out);
  assign zll_main_compute450_in = {zll_main_compute228_in[73:71], zll_main_compute428_out};
  ZLL_Main_compute450  instR4 (zll_main_compute450_in[5:3], zll_main_compute450_in[2:0], zll_main_compute450_out);
  assign resize_inR1 = zll_main_compute450_out;
  assign binop_in = {128'h8, 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h8};
  assign binop_inR3 = {128'(resize_in[63:0]), binop_inR2[255:128] * binop_inR2[127:0]};
  assign resize_inR2 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign zll_main_compute10_in = {zll_main_compute225_in[140:138], zll_main_compute225_in[137:135], zll_main_compute225_in[134:71], zll_main_compute225_in[3:1], zll_main_compute225_in[0]};
  assign resize_inR3 = zll_main_compute10_in[67:4];
  assign zll_main_compute428_inR1 = {zll_main_compute10_in[3:1], zll_main_compute10_in[73:71]};
  ZLL_Main_compute428  instR5 (zll_main_compute428_inR1[5:3], zll_main_compute428_inR1[2:0], zll_main_compute428_outR1);
  assign zll_main_compute450_inR1 = {zll_main_compute10_in[70:68], zll_main_compute428_outR1};
  ZLL_Main_compute450  instR6 (zll_main_compute450_inR1[5:3], zll_main_compute450_inR1[2:0], zll_main_compute450_outR1);
  assign resize_inR4 = zll_main_compute450_outR1;
  assign binop_inR4 = {128'h8, 128'(resize_inR4[2:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h8};
  assign binop_inR7 = {128'(resize_inR3[63:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR5 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign res = (zll_main_compute10_in[0] == 1'h1) ? resize_inR5[7:0] : resize_inR2[7:0];
endmodule

module ZLL_Main_compute119 (input logic [2:0] arg0,
  input logic [63:0] arg1,
  input logic [63:0] arg2,
  input logic [2:0] arg3,
  input logic [2:0] arg4,
  input logic [2:0] arg5,
  output logic [7:0] res);
  logic [5:0] zll_main_compute412_in;
  logic [0:0] zll_main_compute412_out;
  logic [140:0] zll_main_compute364_in;
  logic [5:0] zll_main_compute412_inR1;
  logic [0:0] zll_main_compute412_outR1;
  logic [76:0] zll_main_compute327_in;
  logic [76:0] zll_main_compute384_in;
  logic [63:0] resize_in;
  logic [5:0] zll_main_compute373_in;
  logic [2:0] zll_main_compute373_out;
  logic [5:0] zll_main_compute326_in;
  logic [2:0] zll_main_compute326_out;
  logic [5:0] zll_main_compute450_in;
  logic [2:0] zll_main_compute450_out;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR2;
  logic [73:0] zll_main_compute_in;
  logic [63:0] resize_inR3;
  logic [5:0] zll_main_compute326_inR1;
  logic [2:0] zll_main_compute326_outR1;
  logic [5:0] zll_main_compute450_inR1;
  logic [2:0] zll_main_compute450_outR1;
  logic [2:0] resize_inR4;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR5;
  assign zll_main_compute412_in = {arg5, arg0};
  ZLL_Main_compute412  inst (zll_main_compute412_in[5:3], zll_main_compute412_in[2:0], zll_main_compute412_out);
  assign zll_main_compute364_in = {arg0, arg5, arg1, arg2, arg3, arg4, zll_main_compute412_out};
  assign zll_main_compute412_inR1 = {zll_main_compute364_in[137:135], zll_main_compute364_in[140:138]};
  ZLL_Main_compute412  instR1 (zll_main_compute412_inR1[5:3], zll_main_compute412_inR1[2:0], zll_main_compute412_outR1);
  assign zll_main_compute327_in = {zll_main_compute364_in[140:138], zll_main_compute364_in[137:135], zll_main_compute364_in[134:71], zll_main_compute364_in[6:4], zll_main_compute364_in[3:1], zll_main_compute412_outR1};
  assign zll_main_compute384_in = {zll_main_compute327_in[76:74], zll_main_compute327_in[73:71], zll_main_compute327_in[70:7], zll_main_compute327_in[6:4], zll_main_compute327_in[3:1], zll_main_compute327_in[0]};
  assign resize_in = zll_main_compute384_in[70:7];
  assign zll_main_compute373_in = {zll_main_compute384_in[73:71], zll_main_compute384_in[76:74]};
  ZLL_Main_compute373  instR2 (zll_main_compute373_in[5:3], zll_main_compute373_in[2:0], zll_main_compute373_out);
  assign zll_main_compute326_in = {zll_main_compute373_out, zll_main_compute384_in[3:1]};
  ZLL_Main_compute326  instR3 (zll_main_compute326_in[5:3], zll_main_compute326_in[2:0], zll_main_compute326_out);
  assign zll_main_compute450_in = {zll_main_compute326_out, zll_main_compute384_in[6:4]};
  ZLL_Main_compute450  instR4 (zll_main_compute450_in[5:3], zll_main_compute450_in[2:0], zll_main_compute450_out);
  assign resize_inR1 = zll_main_compute450_out;
  assign binop_in = {128'h8, 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h8};
  assign binop_inR3 = {128'(resize_in[63:0]), binop_inR2[255:128] * binop_inR2[127:0]};
  assign resize_inR2 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign zll_main_compute_in = {zll_main_compute364_in[137:135], zll_main_compute364_in[70:7], zll_main_compute364_in[6:4], zll_main_compute364_in[3:1], zll_main_compute364_in[0]};
  assign resize_inR3 = zll_main_compute_in[70:7];
  assign zll_main_compute326_inR1 = {zll_main_compute_in[73:71], zll_main_compute_in[3:1]};
  ZLL_Main_compute326  instR5 (zll_main_compute326_inR1[5:3], zll_main_compute326_inR1[2:0], zll_main_compute326_outR1);
  assign zll_main_compute450_inR1 = {zll_main_compute326_outR1, zll_main_compute_in[6:4]};
  ZLL_Main_compute450  instR6 (zll_main_compute450_inR1[5:3], zll_main_compute450_inR1[2:0], zll_main_compute450_outR1);
  assign resize_inR4 = zll_main_compute450_outR1;
  assign binop_inR4 = {128'h8, 128'(resize_inR4[2:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h8};
  assign binop_inR7 = {128'(resize_inR3[63:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR5 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign res = (zll_main_compute_in[0] == 1'h1) ? resize_inR5[7:0] : resize_inR2[7:0];
endmodule

module ZLL_Main_compute28 (input logic [63:0] arg0,
  input logic [2:0] arg1,
  input logic [2:0] arg2,
  input logic [2:0] arg3,
  input logic [63:0] arg4,
  input logic [2:0] arg5,
  output logic [7:0] res);
  logic [5:0] zll_main_compute412_in;
  logic [0:0] zll_main_compute412_out;
  logic [140:0] zll_main_compute105_in;
  logic [5:0] zll_main_compute412_inR1;
  logic [0:0] zll_main_compute412_outR1;
  logic [76:0] zll_main_compute431_in;
  logic [76:0] zll_main_compute438_in;
  logic [63:0] resize_in;
  logic [5:0] zll_main_compute373_in;
  logic [2:0] zll_main_compute373_out;
  logic [5:0] zll_main_compute326_in;
  logic [2:0] zll_main_compute326_out;
  logic [5:0] zll_main_compute450_in;
  logic [2:0] zll_main_compute450_out;
  logic [2:0] resize_inR1;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [255:0] binop_inR3;
  logic [127:0] resize_inR2;
  logic [73:0] zll_main_compute222_in;
  logic [63:0] resize_inR3;
  logic [5:0] zll_main_compute326_inR1;
  logic [2:0] zll_main_compute326_outR1;
  logic [5:0] zll_main_compute450_inR1;
  logic [2:0] zll_main_compute450_outR1;
  logic [2:0] resize_inR4;
  logic [255:0] binop_inR4;
  logic [255:0] binop_inR5;
  logic [255:0] binop_inR6;
  logic [255:0] binop_inR7;
  logic [127:0] resize_inR5;
  assign zll_main_compute412_in = {arg5, arg3};
  ZLL_Main_compute412  inst (zll_main_compute412_in[5:3], zll_main_compute412_in[2:0], zll_main_compute412_out);
  assign zll_main_compute105_in = {arg0, arg5, arg1, arg2, arg3, arg4, zll_main_compute412_out};
  assign zll_main_compute412_inR1 = {zll_main_compute105_in[76:74], zll_main_compute105_in[67:65]};
  ZLL_Main_compute412  instR1 (zll_main_compute412_inR1[5:3], zll_main_compute412_inR1[2:0], zll_main_compute412_outR1);
  assign zll_main_compute431_in = {zll_main_compute105_in[140:77], zll_main_compute105_in[76:74], zll_main_compute105_in[73:71], zll_main_compute105_in[70:68], zll_main_compute105_in[67:65], zll_main_compute412_outR1};
  assign zll_main_compute438_in = {zll_main_compute431_in[76:13], zll_main_compute431_in[12:10], zll_main_compute431_in[9:7], zll_main_compute431_in[6:4], zll_main_compute431_in[3:1], zll_main_compute431_in[0]};
  assign resize_in = zll_main_compute438_in[76:13];
  assign zll_main_compute373_in = {zll_main_compute438_in[12:10], zll_main_compute438_in[3:1]};
  ZLL_Main_compute373  instR2 (zll_main_compute373_in[5:3], zll_main_compute373_in[2:0], zll_main_compute373_out);
  assign zll_main_compute326_in = {zll_main_compute373_out, zll_main_compute438_in[6:4]};
  ZLL_Main_compute326  instR3 (zll_main_compute326_in[5:3], zll_main_compute326_in[2:0], zll_main_compute326_out);
  assign zll_main_compute450_in = {zll_main_compute326_out, zll_main_compute438_in[9:7]};
  ZLL_Main_compute450  instR4 (zll_main_compute450_in[5:3], zll_main_compute450_in[2:0], zll_main_compute450_out);
  assign resize_inR1 = zll_main_compute450_out;
  assign binop_in = {128'h8, 128'(resize_inR1[2:0])};
  assign binop_inR1 = {binop_in[255:128] - binop_in[127:0], 128'h1};
  assign binop_inR2 = {binop_inR1[255:128] - binop_inR1[127:0], 128'h8};
  assign binop_inR3 = {128'(resize_in[63:0]), binop_inR2[255:128] * binop_inR2[127:0]};
  assign resize_inR2 = binop_inR3[255:128] >> binop_inR3[127:0];
  assign zll_main_compute222_in = {zll_main_compute105_in[76:74], zll_main_compute105_in[73:71], zll_main_compute105_in[70:68], zll_main_compute105_in[64:1], zll_main_compute105_in[0]};
  assign resize_inR3 = zll_main_compute222_in[64:1];
  assign zll_main_compute326_inR1 = {zll_main_compute222_in[73:71], zll_main_compute222_in[67:65]};
  ZLL_Main_compute326  instR5 (zll_main_compute326_inR1[5:3], zll_main_compute326_inR1[2:0], zll_main_compute326_outR1);
  assign zll_main_compute450_inR1 = {zll_main_compute326_outR1, zll_main_compute222_in[70:68]};
  ZLL_Main_compute450  instR6 (zll_main_compute450_inR1[5:3], zll_main_compute450_inR1[2:0], zll_main_compute450_outR1);
  assign resize_inR4 = zll_main_compute450_outR1;
  assign binop_inR4 = {128'h8, 128'(resize_inR4[2:0])};
  assign binop_inR5 = {binop_inR4[255:128] - binop_inR4[127:0], 128'h1};
  assign binop_inR6 = {binop_inR5[255:128] - binop_inR5[127:0], 128'h8};
  assign binop_inR7 = {128'(resize_inR3[63:0]), binop_inR6[255:128] * binop_inR6[127:0]};
  assign resize_inR5 = binop_inR7[255:128] >> binop_inR7[127:0];
  assign res = (zll_main_compute222_in[0] == 1'h1) ? resize_inR5[7:0] : resize_inR2[7:0];
endmodule