module top_level (input logic [127:0] __in0,
  input logic [127:0] __in1,
  output logic [127:0] __out0);
  logic [255:0] zll_main_multiplyfun1_in;
  logic [255:0] main_multiply_in;
  logic [255:0] zll_main_multiply1304_in;
  logic [255:0] zll_main_multiply1066_in;
  logic [255:0] zll_main_multiply1727_in;
  logic [383:0] zll_main_multiply459_in;
  logic [127:0] id_in;
  logic [384:0] zll_main_multiply1476_in;
  logic [127:0] id_inR1;
  logic [128:0] zll_main_multiply1792_in;
  logic [127:0] zll_main_multiply1792_out;
  logic [256:0] zll_main_multiply1788_in;
  logic [127:0] zll_main_multiply1788_out;
  logic [383:0] zll_main_multiply939_in;
  logic [127:0] id_inR2;
  logic [0:0] rewire_prelude_not_in;
  logic [0:0] rewire_prelude_not_out;
  logic [128:0] zll_main_multiply1785_in;
  logic [127:0] zll_main_multiply1785_out;
  logic [383:0] zll_main_multiply62_in;
  logic [127:0] id_inR3;
  logic [384:0] zll_main_multiply1570_in;
  logic [127:0] id_inR4;
  logic [128:0] zll_main_multiply1792_inR1;
  logic [127:0] zll_main_multiply1792_outR1;
  logic [256:0] zll_main_multiply1749_in;
  logic [127:0] zll_main_multiply1749_out;
  logic [383:0] zll_main_multiply637_in;
  logic [127:0] id_inR5;
  logic [0:0] rewire_prelude_not_inR1;
  logic [0:0] rewire_prelude_not_outR1;
  logic [128:0] zll_main_multiply1785_inR1;
  logic [127:0] zll_main_multiply1785_outR1;
  logic [383:0] zll_main_multiply1342_in;
  logic [127:0] id_inR6;
  logic [384:0] zll_main_multiply811_in;
  logic [127:0] id_inR7;
  logic [128:0] zll_main_multiply1792_inR2;
  logic [127:0] zll_main_multiply1792_outR2;
  logic [256:0] zll_main_multiply1788_inR1;
  logic [127:0] zll_main_multiply1788_outR1;
  logic [383:0] zll_main_multiply681_in;
  logic [127:0] id_inR8;
  logic [0:0] rewire_prelude_not_inR2;
  logic [0:0] rewire_prelude_not_outR2;
  logic [128:0] zll_main_multiply1785_inR2;
  logic [127:0] zll_main_multiply1785_outR2;
  logic [383:0] zll_main_multiply1772_in;
  logic [127:0] id_inR9;
  logic [384:0] zll_main_multiply322_in;
  logic [127:0] id_inR10;
  logic [128:0] zll_main_multiply1792_inR3;
  logic [127:0] zll_main_multiply1792_outR3;
  logic [256:0] zll_main_multiply1788_inR2;
  logic [127:0] zll_main_multiply1788_outR2;
  logic [383:0] zll_main_multiply864_in;
  logic [127:0] id_inR11;
  logic [0:0] rewire_prelude_not_inR3;
  logic [0:0] rewire_prelude_not_outR3;
  logic [128:0] zll_main_multiply1785_inR3;
  logic [127:0] zll_main_multiply1785_outR3;
  logic [383:0] zll_main_multiply516_in;
  logic [127:0] id_inR12;
  logic [384:0] zll_main_multiply1041_in;
  logic [127:0] id_inR13;
  logic [128:0] zll_main_multiply1792_inR4;
  logic [127:0] zll_main_multiply1792_outR4;
  logic [256:0] zll_main_multiply1749_inR1;
  logic [127:0] zll_main_multiply1749_outR1;
  logic [383:0] zll_main_multiply1038_in;
  logic [127:0] id_inR14;
  logic [0:0] rewire_prelude_not_inR4;
  logic [0:0] rewire_prelude_not_outR4;
  logic [128:0] zll_main_multiply1785_inR4;
  logic [127:0] zll_main_multiply1785_outR4;
  logic [383:0] zll_main_multiply151_in;
  logic [127:0] id_inR15;
  logic [384:0] zll_main_multiply909_in;
  logic [127:0] id_inR16;
  logic [128:0] zll_main_multiply1792_inR5;
  logic [127:0] zll_main_multiply1792_outR5;
  logic [256:0] zll_main_multiply1788_inR3;
  logic [127:0] zll_main_multiply1788_outR3;
  logic [383:0] zll_main_multiply1491_in;
  logic [127:0] id_inR17;
  logic [0:0] rewire_prelude_not_inR5;
  logic [0:0] rewire_prelude_not_outR5;
  logic [128:0] zll_main_multiply1785_inR5;
  logic [127:0] zll_main_multiply1785_outR5;
  logic [383:0] zll_main_multiply628_in;
  logic [127:0] id_inR18;
  logic [384:0] zll_main_multiply1395_in;
  logic [127:0] id_inR19;
  logic [128:0] zll_main_multiply1792_inR6;
  logic [127:0] zll_main_multiply1792_outR6;
  logic [256:0] zll_main_multiply1788_inR4;
  logic [127:0] zll_main_multiply1788_outR4;
  logic [383:0] zll_main_multiply305_in;
  logic [127:0] id_inR20;
  logic [0:0] rewire_prelude_not_inR6;
  logic [0:0] rewire_prelude_not_outR6;
  logic [128:0] zll_main_multiply1785_inR6;
  logic [127:0] zll_main_multiply1785_outR6;
  logic [383:0] zll_main_multiply667_in;
  logic [127:0] id_inR21;
  logic [384:0] zll_main_multiply218_in;
  logic [127:0] id_inR22;
  logic [128:0] zll_main_multiply1792_inR7;
  logic [127:0] zll_main_multiply1792_outR7;
  logic [256:0] zll_main_multiply1749_inR2;
  logic [127:0] zll_main_multiply1749_outR2;
  logic [383:0] zll_main_multiply97_in;
  logic [127:0] id_inR23;
  logic [0:0] rewire_prelude_not_inR7;
  logic [0:0] rewire_prelude_not_outR7;
  logic [128:0] zll_main_multiply1785_inR7;
  logic [127:0] zll_main_multiply1785_outR7;
  logic [383:0] zll_main_multiply202_in;
  logic [127:0] id_inR24;
  logic [384:0] zll_main_multiply143_in;
  logic [127:0] id_inR25;
  logic [128:0] zll_main_multiply1792_inR8;
  logic [127:0] zll_main_multiply1792_outR8;
  logic [256:0] zll_main_multiply1788_inR5;
  logic [127:0] zll_main_multiply1788_outR5;
  logic [383:0] zll_main_multiply1630_in;
  logic [127:0] id_inR26;
  logic [0:0] rewire_prelude_not_inR8;
  logic [0:0] rewire_prelude_not_outR8;
  logic [128:0] zll_main_multiply1785_inR8;
  logic [127:0] zll_main_multiply1785_outR8;
  logic [383:0] zll_main_multiply1766_in;
  logic [127:0] id_inR27;
  logic [384:0] zll_main_multiply918_in;
  logic [127:0] id_inR28;
  logic [128:0] zll_main_multiply1792_inR9;
  logic [127:0] zll_main_multiply1792_outR9;
  logic [256:0] zll_main_multiply1788_inR6;
  logic [127:0] zll_main_multiply1788_outR6;
  logic [383:0] zll_main_multiply978_in;
  logic [127:0] id_inR29;
  logic [0:0] rewire_prelude_not_inR9;
  logic [0:0] rewire_prelude_not_outR9;
  logic [128:0] zll_main_multiply1785_inR9;
  logic [127:0] zll_main_multiply1785_outR9;
  logic [383:0] zll_main_multiply497_in;
  logic [127:0] id_inR30;
  logic [384:0] zll_main_multiply617_in;
  logic [127:0] id_inR31;
  logic [128:0] zll_main_multiply1792_inR10;
  logic [127:0] zll_main_multiply1792_outR10;
  logic [256:0] zll_main_multiply1749_inR3;
  logic [127:0] zll_main_multiply1749_outR3;
  logic [383:0] zll_main_multiply1473_in;
  logic [127:0] id_inR32;
  logic [0:0] rewire_prelude_not_inR10;
  logic [0:0] rewire_prelude_not_outR10;
  logic [128:0] zll_main_multiply1785_inR10;
  logic [127:0] zll_main_multiply1785_outR10;
  logic [383:0] zll_main_multiply1206_in;
  logic [127:0] id_inR33;
  logic [384:0] zll_main_multiply158_in;
  logic [127:0] id_inR34;
  logic [128:0] zll_main_multiply1792_inR11;
  logic [127:0] zll_main_multiply1792_outR11;
  logic [256:0] zll_main_multiply1749_inR4;
  logic [127:0] zll_main_multiply1749_outR4;
  logic [383:0] zll_main_multiply769_in;
  logic [127:0] id_inR35;
  logic [0:0] rewire_prelude_not_inR11;
  logic [0:0] rewire_prelude_not_outR11;
  logic [128:0] zll_main_multiply1785_inR11;
  logic [127:0] zll_main_multiply1785_outR11;
  logic [383:0] zll_main_multiply730_in;
  logic [127:0] id_inR36;
  logic [384:0] zll_main_multiply1089_in;
  logic [127:0] id_inR37;
  logic [128:0] zll_main_multiply1792_inR12;
  logic [127:0] zll_main_multiply1792_outR12;
  logic [256:0] zll_main_multiply1749_inR5;
  logic [127:0] zll_main_multiply1749_outR5;
  logic [383:0] zll_main_multiply871_in;
  logic [127:0] id_inR38;
  logic [0:0] rewire_prelude_not_inR12;
  logic [0:0] rewire_prelude_not_outR12;
  logic [128:0] zll_main_multiply1785_inR12;
  logic [127:0] zll_main_multiply1785_outR12;
  logic [383:0] zll_main_multiply279_in;
  logic [127:0] id_inR39;
  logic [384:0] zll_main_multiply39_in;
  logic [127:0] id_inR40;
  logic [128:0] zll_main_multiply1792_inR13;
  logic [127:0] zll_main_multiply1792_outR13;
  logic [256:0] zll_main_multiply1749_inR6;
  logic [127:0] zll_main_multiply1749_outR6;
  logic [383:0] zll_main_multiply1691_in;
  logic [127:0] id_inR41;
  logic [0:0] rewire_prelude_not_inR13;
  logic [0:0] rewire_prelude_not_outR13;
  logic [128:0] zll_main_multiply1785_inR13;
  logic [127:0] zll_main_multiply1785_outR13;
  logic [383:0] zll_main_multiply1282_in;
  logic [127:0] id_inR42;
  logic [384:0] zll_main_multiply110_in;
  logic [127:0] id_inR43;
  logic [128:0] zll_main_multiply1792_inR14;
  logic [127:0] zll_main_multiply1792_outR14;
  logic [256:0] zll_main_multiply1749_inR7;
  logic [127:0] zll_main_multiply1749_outR7;
  logic [383:0] zll_main_multiply282_in;
  logic [127:0] id_inR44;
  logic [0:0] rewire_prelude_not_inR14;
  logic [0:0] rewire_prelude_not_outR14;
  logic [128:0] zll_main_multiply1785_inR14;
  logic [127:0] zll_main_multiply1785_outR14;
  logic [383:0] zll_main_multiply71_in;
  logic [127:0] id_inR45;
  logic [384:0] zll_main_multiply1176_in;
  logic [127:0] id_inR46;
  logic [128:0] zll_main_multiply1792_inR15;
  logic [127:0] zll_main_multiply1792_outR15;
  logic [256:0] zll_main_multiply1788_inR7;
  logic [127:0] zll_main_multiply1788_outR7;
  logic [383:0] zll_main_multiply910_in;
  logic [127:0] id_inR47;
  logic [0:0] rewire_prelude_not_inR15;
  logic [0:0] rewire_prelude_not_outR15;
  logic [128:0] zll_main_multiply1785_inR15;
  logic [127:0] zll_main_multiply1785_outR15;
  logic [383:0] zll_main_multiply1165_in;
  logic [127:0] id_inR48;
  logic [384:0] zll_main_multiply168_in;
  logic [127:0] id_inR49;
  logic [128:0] zll_main_multiply1792_inR16;
  logic [127:0] zll_main_multiply1792_outR16;
  logic [256:0] zll_main_multiply1788_inR8;
  logic [127:0] zll_main_multiply1788_outR8;
  logic [383:0] zll_main_multiply195_in;
  logic [127:0] id_inR50;
  logic [0:0] rewire_prelude_not_inR16;
  logic [0:0] rewire_prelude_not_outR16;
  logic [128:0] zll_main_multiply1785_inR16;
  logic [127:0] zll_main_multiply1785_outR16;
  logic [383:0] zll_main_multiply750_in;
  logic [127:0] id_inR51;
  logic [384:0] zll_main_multiply196_in;
  logic [127:0] id_inR52;
  logic [128:0] zll_main_multiply1792_inR17;
  logic [127:0] zll_main_multiply1792_outR17;
  logic [256:0] zll_main_multiply1788_inR9;
  logic [127:0] zll_main_multiply1788_outR9;
  logic [383:0] zll_main_multiply765_in;
  logic [127:0] id_inR53;
  logic [0:0] rewire_prelude_not_inR17;
  logic [0:0] rewire_prelude_not_outR17;
  logic [128:0] zll_main_multiply1785_inR17;
  logic [127:0] zll_main_multiply1785_outR17;
  logic [383:0] zll_main_multiply851_in;
  logic [127:0] id_inR54;
  logic [384:0] zll_main_multiply831_in;
  logic [127:0] id_inR55;
  logic [128:0] zll_main_multiply1792_inR18;
  logic [127:0] zll_main_multiply1792_outR18;
  logic [256:0] zll_main_multiply1788_inR10;
  logic [127:0] zll_main_multiply1788_outR10;
  logic [383:0] zll_main_multiply1107_in;
  logic [127:0] id_inR56;
  logic [0:0] rewire_prelude_not_inR18;
  logic [0:0] rewire_prelude_not_outR18;
  logic [128:0] zll_main_multiply1785_inR18;
  logic [127:0] zll_main_multiply1785_outR18;
  logic [383:0] zll_main_multiply29_in;
  logic [127:0] id_inR57;
  logic [384:0] zll_main_multiply964_in;
  logic [127:0] id_inR58;
  logic [128:0] zll_main_multiply1792_inR19;
  logic [127:0] zll_main_multiply1792_outR19;
  logic [256:0] zll_main_multiply1788_inR11;
  logic [127:0] zll_main_multiply1788_outR11;
  logic [383:0] zll_main_multiply1345_in;
  logic [127:0] id_inR59;
  logic [0:0] rewire_prelude_not_inR19;
  logic [0:0] rewire_prelude_not_outR19;
  logic [128:0] zll_main_multiply1785_inR19;
  logic [127:0] zll_main_multiply1785_outR19;
  logic [383:0] zll_main_multiply390_in;
  logic [127:0] id_inR60;
  logic [384:0] zll_main_multiply1076_in;
  logic [127:0] id_inR61;
  logic [128:0] zll_main_multiply1792_inR20;
  logic [127:0] zll_main_multiply1792_outR20;
  logic [256:0] zll_main_multiply1749_inR8;
  logic [127:0] zll_main_multiply1749_outR8;
  logic [383:0] zll_main_multiply687_in;
  logic [127:0] id_inR62;
  logic [0:0] rewire_prelude_not_inR20;
  logic [0:0] rewire_prelude_not_outR20;
  logic [128:0] zll_main_multiply1785_inR20;
  logic [127:0] zll_main_multiply1785_outR20;
  logic [383:0] zll_main_multiply138_in;
  logic [127:0] id_inR63;
  logic [384:0] zll_main_multiply1411_in;
  logic [127:0] id_inR64;
  logic [128:0] zll_main_multiply1792_inR21;
  logic [127:0] zll_main_multiply1792_outR21;
  logic [256:0] zll_main_multiply1788_inR12;
  logic [127:0] zll_main_multiply1788_outR12;
  logic [383:0] zll_main_multiply101_in;
  logic [127:0] id_inR65;
  logic [0:0] rewire_prelude_not_inR21;
  logic [0:0] rewire_prelude_not_outR21;
  logic [128:0] zll_main_multiply1785_inR21;
  logic [127:0] zll_main_multiply1785_outR21;
  logic [383:0] zll_main_multiply686_in;
  logic [127:0] id_inR66;
  logic [384:0] zll_main_multiply1013_in;
  logic [127:0] id_inR67;
  logic [128:0] zll_main_multiply1792_inR22;
  logic [127:0] zll_main_multiply1792_outR22;
  logic [256:0] zll_main_multiply1788_inR13;
  logic [127:0] zll_main_multiply1788_outR13;
  logic [383:0] zll_main_multiply1487_in;
  logic [127:0] id_inR68;
  logic [0:0] rewire_prelude_not_inR22;
  logic [0:0] rewire_prelude_not_outR22;
  logic [128:0] zll_main_multiply1785_inR22;
  logic [127:0] zll_main_multiply1785_outR22;
  logic [383:0] zll_main_multiply178_in;
  logic [127:0] id_inR69;
  logic [384:0] zll_main_multiply952_in;
  logic [127:0] id_inR70;
  logic [128:0] zll_main_multiply1792_inR23;
  logic [127:0] zll_main_multiply1792_outR23;
  logic [256:0] zll_main_multiply1749_inR9;
  logic [127:0] zll_main_multiply1749_outR9;
  logic [383:0] zll_main_multiply148_in;
  logic [127:0] id_inR71;
  logic [0:0] rewire_prelude_not_inR23;
  logic [0:0] rewire_prelude_not_outR23;
  logic [128:0] zll_main_multiply1785_inR23;
  logic [127:0] zll_main_multiply1785_outR23;
  logic [383:0] zll_main_multiply485_in;
  logic [127:0] id_inR72;
  logic [384:0] zll_main_multiply1592_in;
  logic [127:0] id_inR73;
  logic [128:0] zll_main_multiply1792_inR24;
  logic [127:0] zll_main_multiply1792_outR24;
  logic [256:0] zll_main_multiply1788_inR14;
  logic [127:0] zll_main_multiply1788_outR14;
  logic [383:0] zll_main_multiply879_in;
  logic [127:0] id_inR74;
  logic [0:0] rewire_prelude_not_inR24;
  logic [0:0] rewire_prelude_not_outR24;
  logic [128:0] zll_main_multiply1785_inR24;
  logic [127:0] zll_main_multiply1785_outR24;
  logic [383:0] zll_main_multiply1327_in;
  logic [127:0] id_inR75;
  logic [384:0] zll_main_multiply724_in;
  logic [127:0] id_inR76;
  logic [128:0] zll_main_multiply1792_inR25;
  logic [127:0] zll_main_multiply1792_outR25;
  logic [256:0] zll_main_multiply1749_inR10;
  logic [127:0] zll_main_multiply1749_outR10;
  logic [383:0] zll_main_multiply904_in;
  logic [127:0] id_inR77;
  logic [0:0] rewire_prelude_not_inR25;
  logic [0:0] rewire_prelude_not_outR25;
  logic [128:0] zll_main_multiply1785_inR25;
  logic [127:0] zll_main_multiply1785_outR25;
  logic [383:0] zll_main_multiply705_in;
  logic [127:0] id_inR78;
  logic [384:0] zll_main_multiply627_in;
  logic [127:0] id_inR79;
  logic [128:0] zll_main_multiply1792_inR26;
  logic [127:0] zll_main_multiply1792_outR26;
  logic [256:0] zll_main_multiply1788_inR15;
  logic [127:0] zll_main_multiply1788_outR15;
  logic [383:0] zll_main_multiply847_in;
  logic [127:0] id_inR80;
  logic [0:0] rewire_prelude_not_inR26;
  logic [0:0] rewire_prelude_not_outR26;
  logic [128:0] zll_main_multiply1785_inR26;
  logic [127:0] zll_main_multiply1785_outR26;
  logic [383:0] zll_main_multiply560_in;
  logic [127:0] id_inR81;
  logic [384:0] zll_main_multiply901_in;
  logic [127:0] id_inR82;
  logic [128:0] zll_main_multiply1792_inR27;
  logic [127:0] zll_main_multiply1792_outR27;
  logic [256:0] zll_main_multiply1788_inR16;
  logic [127:0] zll_main_multiply1788_outR16;
  logic [383:0] zll_main_multiply420_in;
  logic [127:0] id_inR83;
  logic [0:0] rewire_prelude_not_inR27;
  logic [0:0] rewire_prelude_not_outR27;
  logic [128:0] zll_main_multiply1785_inR27;
  logic [127:0] zll_main_multiply1785_outR27;
  logic [383:0] zll_main_multiply291_in;
  logic [127:0] id_inR84;
  logic [384:0] zll_main_multiply185_in;
  logic [127:0] id_inR85;
  logic [128:0] zll_main_multiply1792_inR28;
  logic [127:0] zll_main_multiply1792_outR28;
  logic [256:0] zll_main_multiply1788_inR17;
  logic [127:0] zll_main_multiply1788_outR17;
  logic [383:0] zll_main_multiply749_in;
  logic [127:0] id_inR86;
  logic [0:0] rewire_prelude_not_inR28;
  logic [0:0] rewire_prelude_not_outR28;
  logic [128:0] zll_main_multiply1785_inR28;
  logic [127:0] zll_main_multiply1785_outR28;
  logic [383:0] zll_main_multiply810_in;
  logic [127:0] id_inR87;
  logic [384:0] zll_main_multiply154_in;
  logic [127:0] id_inR88;
  logic [128:0] zll_main_multiply1792_inR29;
  logic [127:0] zll_main_multiply1792_outR29;
  logic [256:0] zll_main_multiply1749_inR11;
  logic [127:0] zll_main_multiply1749_outR11;
  logic [383:0] zll_main_multiply1542_in;
  logic [127:0] id_inR89;
  logic [0:0] rewire_prelude_not_inR29;
  logic [0:0] rewire_prelude_not_outR29;
  logic [128:0] zll_main_multiply1785_inR29;
  logic [127:0] zll_main_multiply1785_outR29;
  logic [383:0] zll_main_multiply1173_in;
  logic [127:0] id_inR90;
  logic [384:0] zll_main_multiply512_in;
  logic [127:0] id_inR91;
  logic [128:0] zll_main_multiply1792_inR30;
  logic [127:0] zll_main_multiply1792_outR30;
  logic [256:0] zll_main_multiply1788_inR18;
  logic [127:0] zll_main_multiply1788_outR18;
  logic [383:0] zll_main_multiply66_in;
  logic [127:0] id_inR92;
  logic [0:0] rewire_prelude_not_inR30;
  logic [0:0] rewire_prelude_not_outR30;
  logic [128:0] zll_main_multiply1785_inR30;
  logic [127:0] zll_main_multiply1785_outR30;
  logic [383:0] zll_main_multiply1574_in;
  logic [127:0] id_inR93;
  logic [384:0] zll_main_multiply550_in;
  logic [127:0] id_inR94;
  logic [128:0] zll_main_multiply1792_inR31;
  logic [127:0] zll_main_multiply1792_outR31;
  logic [256:0] zll_main_multiply1788_inR19;
  logic [127:0] zll_main_multiply1788_outR19;
  logic [383:0] zll_main_multiply1392_in;
  logic [127:0] id_inR95;
  logic [0:0] rewire_prelude_not_inR31;
  logic [0:0] rewire_prelude_not_outR31;
  logic [128:0] zll_main_multiply1785_inR31;
  logic [127:0] zll_main_multiply1785_outR31;
  logic [383:0] zll_main_multiply450_in;
  logic [127:0] id_inR96;
  logic [384:0] zll_main_multiply193_in;
  logic [127:0] id_inR97;
  logic [128:0] zll_main_multiply1792_inR32;
  logic [127:0] zll_main_multiply1792_outR32;
  logic [256:0] zll_main_multiply1788_inR20;
  logic [127:0] zll_main_multiply1788_outR20;
  logic [383:0] zll_main_multiply633_in;
  logic [127:0] id_inR98;
  logic [0:0] rewire_prelude_not_inR32;
  logic [0:0] rewire_prelude_not_outR32;
  logic [128:0] zll_main_multiply1785_inR32;
  logic [127:0] zll_main_multiply1785_outR32;
  logic [383:0] zll_main_multiply1596_in;
  logic [127:0] id_inR99;
  logic [384:0] zll_main_multiply315_in;
  logic [127:0] id_inR100;
  logic [128:0] zll_main_multiply1792_inR33;
  logic [127:0] zll_main_multiply1792_outR33;
  logic [256:0] zll_main_multiply1749_inR12;
  logic [127:0] zll_main_multiply1749_outR12;
  logic [383:0] zll_main_multiply165_in;
  logic [127:0] id_inR101;
  logic [0:0] rewire_prelude_not_inR33;
  logic [0:0] rewire_prelude_not_outR33;
  logic [128:0] zll_main_multiply1785_inR33;
  logic [127:0] zll_main_multiply1785_outR33;
  logic [383:0] zll_main_multiply934_in;
  logic [127:0] id_inR102;
  logic [384:0] zll_main_multiply738_in;
  logic [127:0] id_inR103;
  logic [128:0] zll_main_multiply1792_inR34;
  logic [127:0] zll_main_multiply1792_outR34;
  logic [256:0] zll_main_multiply1788_inR21;
  logic [127:0] zll_main_multiply1788_outR21;
  logic [383:0] zll_main_multiply278_in;
  logic [127:0] id_inR104;
  logic [0:0] rewire_prelude_not_inR34;
  logic [0:0] rewire_prelude_not_outR34;
  logic [128:0] zll_main_multiply1785_inR34;
  logic [127:0] zll_main_multiply1785_outR34;
  logic [383:0] zll_main_multiply271_in;
  logic [127:0] id_inR105;
  logic [384:0] zll_main_multiply1331_in;
  logic [127:0] id_inR106;
  logic [128:0] zll_main_multiply1792_inR35;
  logic [127:0] zll_main_multiply1792_outR35;
  logic [256:0] zll_main_multiply1788_inR22;
  logic [127:0] zll_main_multiply1788_outR22;
  logic [383:0] zll_main_multiply993_in;
  logic [127:0] id_inR107;
  logic [0:0] rewire_prelude_not_inR35;
  logic [0:0] rewire_prelude_not_outR35;
  logic [128:0] zll_main_multiply1785_inR35;
  logic [127:0] zll_main_multiply1785_outR35;
  logic [383:0] zll_main_multiply1389_in;
  logic [127:0] id_inR108;
  logic [384:0] zll_main_multiply1343_in;
  logic [127:0] id_inR109;
  logic [128:0] zll_main_multiply1792_inR36;
  logic [127:0] zll_main_multiply1792_outR36;
  logic [256:0] zll_main_multiply1749_inR13;
  logic [127:0] zll_main_multiply1749_outR13;
  logic [383:0] zll_main_multiply873_in;
  logic [127:0] id_inR110;
  logic [0:0] rewire_prelude_not_inR36;
  logic [0:0] rewire_prelude_not_outR36;
  logic [128:0] zll_main_multiply1785_inR36;
  logic [127:0] zll_main_multiply1785_outR36;
  logic [383:0] zll_main_multiply1626_in;
  logic [127:0] id_inR111;
  logic [384:0] zll_main_multiply350_in;
  logic [127:0] id_inR112;
  logic [128:0] zll_main_multiply1792_inR37;
  logic [127:0] zll_main_multiply1792_outR37;
  logic [256:0] zll_main_multiply1749_inR14;
  logic [127:0] zll_main_multiply1749_outR14;
  logic [383:0] zll_main_multiply421_in;
  logic [127:0] id_inR113;
  logic [0:0] rewire_prelude_not_inR37;
  logic [0:0] rewire_prelude_not_outR37;
  logic [128:0] zll_main_multiply1785_inR37;
  logic [127:0] zll_main_multiply1785_outR37;
  logic [383:0] zll_main_multiply556_in;
  logic [127:0] id_inR114;
  logic [384:0] zll_main_multiply1036_in;
  logic [127:0] id_inR115;
  logic [128:0] zll_main_multiply1792_inR38;
  logic [127:0] zll_main_multiply1792_outR38;
  logic [256:0] zll_main_multiply1749_inR15;
  logic [127:0] zll_main_multiply1749_outR15;
  logic [383:0] zll_main_multiply22_in;
  logic [127:0] id_inR116;
  logic [0:0] rewire_prelude_not_inR38;
  logic [0:0] rewire_prelude_not_outR38;
  logic [128:0] zll_main_multiply1785_inR38;
  logic [127:0] zll_main_multiply1785_outR38;
  logic [383:0] zll_main_multiply905_in;
  logic [127:0] id_inR117;
  logic [384:0] zll_main_multiply1518_in;
  logic [127:0] id_inR118;
  logic [128:0] zll_main_multiply1792_inR39;
  logic [127:0] zll_main_multiply1792_outR39;
  logic [256:0] zll_main_multiply1749_inR16;
  logic [127:0] zll_main_multiply1749_outR16;
  logic [383:0] zll_main_multiply403_in;
  logic [127:0] id_inR119;
  logic [0:0] rewire_prelude_not_inR39;
  logic [0:0] rewire_prelude_not_outR39;
  logic [128:0] zll_main_multiply1785_inR39;
  logic [127:0] zll_main_multiply1785_outR39;
  logic [383:0] zll_main_multiply644_in;
  logic [127:0] id_inR120;
  logic [384:0] zll_main_multiply431_in;
  logic [127:0] id_inR121;
  logic [128:0] zll_main_multiply1792_inR40;
  logic [127:0] zll_main_multiply1792_outR40;
  logic [256:0] zll_main_multiply1749_inR17;
  logic [127:0] zll_main_multiply1749_outR17;
  logic [383:0] zll_main_multiply256_in;
  logic [127:0] id_inR122;
  logic [0:0] rewire_prelude_not_inR40;
  logic [0:0] rewire_prelude_not_outR40;
  logic [128:0] zll_main_multiply1785_inR40;
  logic [127:0] zll_main_multiply1785_outR40;
  logic [383:0] zll_main_multiply198_in;
  logic [127:0] id_inR123;
  logic [384:0] zll_main_multiply846_in;
  logic [127:0] id_inR124;
  logic [128:0] zll_main_multiply1792_inR41;
  logic [127:0] zll_main_multiply1792_outR41;
  logic [256:0] zll_main_multiply1749_inR18;
  logic [127:0] zll_main_multiply1749_outR18;
  logic [383:0] zll_main_multiply25_in;
  logic [127:0] id_inR125;
  logic [0:0] rewire_prelude_not_inR41;
  logic [0:0] rewire_prelude_not_outR41;
  logic [128:0] zll_main_multiply1785_inR41;
  logic [127:0] zll_main_multiply1785_outR41;
  logic [383:0] zll_main_multiply381_in;
  logic [127:0] id_inR126;
  logic [384:0] zll_main_multiply285_in;
  logic [127:0] id_inR127;
  logic [128:0] zll_main_multiply1792_inR42;
  logic [127:0] zll_main_multiply1792_outR42;
  logic [256:0] zll_main_multiply1788_inR23;
  logic [127:0] zll_main_multiply1788_outR23;
  logic [383:0] zll_main_multiply1355_in;
  logic [127:0] id_inR128;
  logic [0:0] rewire_prelude_not_inR42;
  logic [0:0] rewire_prelude_not_outR42;
  logic [128:0] zll_main_multiply1785_inR42;
  logic [127:0] zll_main_multiply1785_outR42;
  logic [383:0] zll_main_multiply1141_in;
  logic [127:0] id_inR129;
  logic [384:0] zll_main_multiply188_in;
  logic [127:0] id_inR130;
  logic [128:0] zll_main_multiply1792_inR43;
  logic [127:0] zll_main_multiply1792_outR43;
  logic [256:0] zll_main_multiply1788_inR24;
  logic [127:0] zll_main_multiply1788_outR24;
  logic [383:0] zll_main_multiply558_in;
  logic [127:0] id_inR131;
  logic [0:0] rewire_prelude_not_inR43;
  logic [0:0] rewire_prelude_not_outR43;
  logic [128:0] zll_main_multiply1785_inR43;
  logic [127:0] zll_main_multiply1785_outR43;
  logic [383:0] zll_main_multiply706_in;
  logic [127:0] id_inR132;
  logic [384:0] zll_main_multiply323_in;
  logic [127:0] id_inR133;
  logic [128:0] zll_main_multiply1792_inR44;
  logic [127:0] zll_main_multiply1792_outR44;
  logic [256:0] zll_main_multiply1749_inR19;
  logic [127:0] zll_main_multiply1749_outR19;
  logic [383:0] zll_main_multiply1675_in;
  logic [127:0] id_inR134;
  logic [0:0] rewire_prelude_not_inR44;
  logic [0:0] rewire_prelude_not_outR44;
  logic [128:0] zll_main_multiply1785_inR44;
  logic [127:0] zll_main_multiply1785_outR44;
  logic [383:0] zll_main_multiply863_in;
  logic [127:0] id_inR135;
  logic [384:0] zll_main_multiply1246_in;
  logic [127:0] id_inR136;
  logic [128:0] zll_main_multiply1792_inR45;
  logic [127:0] zll_main_multiply1792_outR45;
  logic [256:0] zll_main_multiply1749_inR20;
  logic [127:0] zll_main_multiply1749_outR20;
  logic [383:0] zll_main_multiply190_in;
  logic [127:0] id_inR137;
  logic [0:0] rewire_prelude_not_inR45;
  logic [0:0] rewire_prelude_not_outR45;
  logic [128:0] zll_main_multiply1785_inR45;
  logic [127:0] zll_main_multiply1785_outR45;
  logic [383:0] zll_main_multiply7_in;
  logic [127:0] id_inR138;
  logic [384:0] zll_main_multiply1112_in;
  logic [127:0] id_inR139;
  logic [128:0] zll_main_multiply1792_inR46;
  logic [127:0] zll_main_multiply1792_outR46;
  logic [256:0] zll_main_multiply1749_inR21;
  logic [127:0] zll_main_multiply1749_outR21;
  logic [383:0] zll_main_multiply906_in;
  logic [127:0] id_inR140;
  logic [0:0] rewire_prelude_not_inR46;
  logic [0:0] rewire_prelude_not_outR46;
  logic [128:0] zll_main_multiply1785_inR46;
  logic [127:0] zll_main_multiply1785_outR46;
  logic [383:0] zll_main_multiply865_in;
  logic [127:0] id_inR141;
  logic [384:0] zll_main_multiply1034_in;
  logic [127:0] id_inR142;
  logic [128:0] zll_main_multiply1792_inR47;
  logic [127:0] zll_main_multiply1792_outR47;
  logic [256:0] zll_main_multiply1788_inR25;
  logic [127:0] zll_main_multiply1788_outR25;
  logic [383:0] zll_main_multiply1238_in;
  logic [127:0] id_inR143;
  logic [0:0] rewire_prelude_not_inR47;
  logic [0:0] rewire_prelude_not_outR47;
  logic [128:0] zll_main_multiply1785_inR47;
  logic [127:0] zll_main_multiply1785_outR47;
  logic [383:0] zll_main_multiply1103_in;
  logic [127:0] id_inR144;
  logic [384:0] zll_main_multiply413_in;
  logic [127:0] id_inR145;
  logic [128:0] zll_main_multiply1792_inR48;
  logic [127:0] zll_main_multiply1792_outR48;
  logic [256:0] zll_main_multiply1749_inR22;
  logic [127:0] zll_main_multiply1749_outR22;
  logic [383:0] zll_main_multiply1177_in;
  logic [127:0] id_inR146;
  logic [0:0] rewire_prelude_not_inR48;
  logic [0:0] rewire_prelude_not_outR48;
  logic [128:0] zll_main_multiply1785_inR48;
  logic [127:0] zll_main_multiply1785_outR48;
  logic [383:0] zll_main_multiply716_in;
  logic [127:0] id_inR147;
  logic [384:0] zll_main_multiply384_in;
  logic [127:0] id_inR148;
  logic [128:0] zll_main_multiply1792_inR49;
  logic [127:0] zll_main_multiply1792_outR49;
  logic [256:0] zll_main_multiply1749_inR23;
  logic [127:0] zll_main_multiply1749_outR23;
  logic [383:0] zll_main_multiply267_in;
  logic [127:0] id_inR149;
  logic [0:0] rewire_prelude_not_inR49;
  logic [0:0] rewire_prelude_not_outR49;
  logic [128:0] zll_main_multiply1785_inR49;
  logic [127:0] zll_main_multiply1785_outR49;
  logic [383:0] zll_main_multiply72_in;
  logic [127:0] id_inR150;
  logic [384:0] zll_main_multiply928_in;
  logic [127:0] id_inR151;
  logic [128:0] zll_main_multiply1792_inR50;
  logic [127:0] zll_main_multiply1792_outR50;
  logic [256:0] zll_main_multiply1788_inR26;
  logic [127:0] zll_main_multiply1788_outR26;
  logic [383:0] zll_main_multiply849_in;
  logic [127:0] id_inR152;
  logic [0:0] rewire_prelude_not_inR50;
  logic [0:0] rewire_prelude_not_outR50;
  logic [128:0] zll_main_multiply1785_inR50;
  logic [127:0] zll_main_multiply1785_outR50;
  logic [383:0] zll_main_multiply1488_in;
  logic [127:0] id_inR153;
  logic [384:0] zll_main_multiply996_in;
  logic [127:0] id_inR154;
  logic [128:0] zll_main_multiply1792_inR51;
  logic [127:0] zll_main_multiply1792_outR51;
  logic [256:0] zll_main_multiply1749_inR24;
  logic [127:0] zll_main_multiply1749_outR24;
  logic [383:0] zll_main_multiply287_in;
  logic [127:0] id_inR155;
  logic [0:0] rewire_prelude_not_inR51;
  logic [0:0] rewire_prelude_not_outR51;
  logic [128:0] zll_main_multiply1785_inR51;
  logic [127:0] zll_main_multiply1785_outR51;
  logic [383:0] zll_main_multiply1648_in;
  logic [127:0] id_inR156;
  logic [384:0] zll_main_multiply868_in;
  logic [127:0] id_inR157;
  logic [128:0] zll_main_multiply1792_inR52;
  logic [127:0] zll_main_multiply1792_outR52;
  logic [256:0] zll_main_multiply1749_inR25;
  logic [127:0] zll_main_multiply1749_outR25;
  logic [383:0] zll_main_multiply594_in;
  logic [127:0] id_inR158;
  logic [0:0] rewire_prelude_not_inR52;
  logic [0:0] rewire_prelude_not_outR52;
  logic [128:0] zll_main_multiply1785_inR52;
  logic [127:0] zll_main_multiply1785_outR52;
  logic [383:0] zll_main_multiply1745_in;
  logic [127:0] id_inR159;
  logic [384:0] zll_main_multiply976_in;
  logic [127:0] id_inR160;
  logic [128:0] zll_main_multiply1792_inR53;
  logic [127:0] zll_main_multiply1792_outR53;
  logic [256:0] zll_main_multiply1788_inR27;
  logic [127:0] zll_main_multiply1788_outR27;
  logic [383:0] zll_main_multiply436_in;
  logic [127:0] id_inR161;
  logic [0:0] rewire_prelude_not_inR53;
  logic [0:0] rewire_prelude_not_outR53;
  logic [128:0] zll_main_multiply1785_inR53;
  logic [127:0] zll_main_multiply1785_outR53;
  logic [383:0] zll_main_multiply260_in;
  logic [127:0] id_inR162;
  logic [384:0] zll_main_multiply1381_in;
  logic [127:0] id_inR163;
  logic [128:0] zll_main_multiply1792_inR54;
  logic [127:0] zll_main_multiply1792_outR54;
  logic [256:0] zll_main_multiply1788_inR28;
  logic [127:0] zll_main_multiply1788_outR28;
  logic [383:0] zll_main_multiply1598_in;
  logic [127:0] id_inR164;
  logic [0:0] rewire_prelude_not_inR54;
  logic [0:0] rewire_prelude_not_outR54;
  logic [128:0] zll_main_multiply1785_inR54;
  logic [127:0] zll_main_multiply1785_outR54;
  logic [383:0] zll_main_multiply1610_in;
  logic [127:0] id_inR165;
  logic [384:0] zll_main_multiply806_in;
  logic [127:0] id_inR166;
  logic [128:0] zll_main_multiply1792_inR55;
  logic [127:0] zll_main_multiply1792_outR55;
  logic [256:0] zll_main_multiply1788_inR29;
  logic [127:0] zll_main_multiply1788_outR29;
  logic [383:0] zll_main_multiply830_in;
  logic [127:0] id_inR167;
  logic [0:0] rewire_prelude_not_inR55;
  logic [0:0] rewire_prelude_not_outR55;
  logic [128:0] zll_main_multiply1785_inR55;
  logic [127:0] zll_main_multiply1785_outR55;
  logic [383:0] zll_main_multiply792_in;
  logic [127:0] id_inR168;
  logic [384:0] zll_main_multiply1584_in;
  logic [127:0] id_inR169;
  logic [128:0] zll_main_multiply1792_inR56;
  logic [127:0] zll_main_multiply1792_outR56;
  logic [256:0] zll_main_multiply1749_inR26;
  logic [127:0] zll_main_multiply1749_outR26;
  logic [383:0] zll_main_multiply14_in;
  logic [127:0] id_inR170;
  logic [0:0] rewire_prelude_not_inR56;
  logic [0:0] rewire_prelude_not_outR56;
  logic [128:0] zll_main_multiply1785_inR56;
  logic [127:0] zll_main_multiply1785_outR56;
  logic [383:0] zll_main_multiply1099_in;
  logic [127:0] id_inR171;
  logic [384:0] zll_main_multiply719_in;
  logic [127:0] id_inR172;
  logic [128:0] zll_main_multiply1792_inR57;
  logic [127:0] zll_main_multiply1792_outR57;
  logic [256:0] zll_main_multiply1749_inR27;
  logic [127:0] zll_main_multiply1749_outR27;
  logic [383:0] zll_main_multiply150_in;
  logic [127:0] id_inR173;
  logic [0:0] rewire_prelude_not_inR57;
  logic [0:0] rewire_prelude_not_outR57;
  logic [128:0] zll_main_multiply1785_inR57;
  logic [127:0] zll_main_multiply1785_outR57;
  logic [383:0] zll_main_multiply1791_in;
  logic [127:0] id_inR174;
  logic [384:0] zll_main_multiply472_in;
  logic [127:0] id_inR175;
  logic [128:0] zll_main_multiply1792_inR58;
  logic [127:0] zll_main_multiply1792_outR58;
  logic [256:0] zll_main_multiply1749_inR28;
  logic [127:0] zll_main_multiply1749_outR28;
  logic [383:0] zll_main_multiply1270_in;
  logic [127:0] id_inR176;
  logic [0:0] rewire_prelude_not_inR58;
  logic [0:0] rewire_prelude_not_outR58;
  logic [128:0] zll_main_multiply1785_inR58;
  logic [127:0] zll_main_multiply1785_outR58;
  logic [383:0] zll_main_multiply1207_in;
  logic [127:0] id_inR177;
  logic [384:0] zll_main_multiply1210_in;
  logic [127:0] id_inR178;
  logic [128:0] zll_main_multiply1792_inR59;
  logic [127:0] zll_main_multiply1792_outR59;
  logic [256:0] zll_main_multiply1788_inR30;
  logic [127:0] zll_main_multiply1788_outR30;
  logic [383:0] zll_main_multiply215_in;
  logic [127:0] id_inR179;
  logic [0:0] rewire_prelude_not_inR59;
  logic [0:0] rewire_prelude_not_outR59;
  logic [128:0] zll_main_multiply1785_inR59;
  logic [127:0] zll_main_multiply1785_outR59;
  logic [383:0] zll_main_multiply1202_in;
  logic [127:0] id_inR180;
  logic [384:0] zll_main_multiply28_in;
  logic [127:0] id_inR181;
  logic [128:0] zll_main_multiply1792_inR60;
  logic [127:0] zll_main_multiply1792_outR60;
  logic [256:0] zll_main_multiply1749_inR29;
  logic [127:0] zll_main_multiply1749_outR29;
  logic [383:0] zll_main_multiply9_in;
  logic [127:0] id_inR182;
  logic [0:0] rewire_prelude_not_inR60;
  logic [0:0] rewire_prelude_not_outR60;
  logic [128:0] zll_main_multiply1785_inR60;
  logic [127:0] zll_main_multiply1785_outR60;
  logic [383:0] zll_main_multiply1279_in;
  logic [127:0] id_inR183;
  logic [384:0] zll_main_multiply132_in;
  logic [127:0] id_inR184;
  logic [128:0] zll_main_multiply1792_inR61;
  logic [127:0] zll_main_multiply1792_outR61;
  logic [256:0] zll_main_multiply1749_inR30;
  logic [127:0] zll_main_multiply1749_outR30;
  logic [383:0] zll_main_multiply530_in;
  logic [127:0] id_inR185;
  logic [0:0] rewire_prelude_not_inR61;
  logic [0:0] rewire_prelude_not_outR61;
  logic [128:0] zll_main_multiply1785_inR61;
  logic [127:0] zll_main_multiply1785_outR61;
  logic [383:0] zll_main_multiply1445_in;
  logic [127:0] id_inR186;
  logic [384:0] zll_main_multiply1545_in;
  logic [127:0] id_inR187;
  logic [128:0] zll_main_multiply1792_inR62;
  logic [127:0] zll_main_multiply1792_outR62;
  logic [256:0] zll_main_multiply1788_inR31;
  logic [127:0] zll_main_multiply1788_outR31;
  logic [383:0] zll_main_multiply1517_in;
  logic [127:0] id_inR188;
  logic [0:0] rewire_prelude_not_inR62;
  logic [0:0] rewire_prelude_not_outR62;
  logic [128:0] zll_main_multiply1785_inR62;
  logic [127:0] zll_main_multiply1785_outR62;
  logic [383:0] zll_main_multiply326_in;
  logic [127:0] id_inR189;
  logic [384:0] zll_main_multiply1468_in;
  logic [127:0] id_inR190;
  logic [128:0] zll_main_multiply1792_inR63;
  logic [127:0] zll_main_multiply1792_outR63;
  logic [256:0] zll_main_multiply1788_inR32;
  logic [127:0] zll_main_multiply1788_outR32;
  logic [383:0] zll_main_multiply1693_in;
  logic [127:0] id_inR191;
  logic [0:0] rewire_prelude_not_inR63;
  logic [0:0] rewire_prelude_not_outR63;
  logic [128:0] zll_main_multiply1785_inR63;
  logic [127:0] zll_main_multiply1785_outR63;
  logic [383:0] zll_main_multiply284_in;
  logic [127:0] id_inR192;
  logic [384:0] zll_main_multiply1639_in;
  logic [127:0] id_inR193;
  logic [128:0] zll_main_multiply1792_inR64;
  logic [127:0] zll_main_multiply1792_outR64;
  logic [256:0] zll_main_multiply1788_inR33;
  logic [127:0] zll_main_multiply1788_outR33;
  logic [383:0] zll_main_multiply675_in;
  logic [127:0] id_inR194;
  logic [0:0] rewire_prelude_not_inR64;
  logic [0:0] rewire_prelude_not_outR64;
  logic [128:0] zll_main_multiply1785_inR64;
  logic [127:0] zll_main_multiply1785_outR64;
  logic [383:0] zll_main_multiply1633_in;
  logic [127:0] id_inR195;
  logic [384:0] zll_main_multiply1469_in;
  logic [127:0] id_inR196;
  logic [128:0] zll_main_multiply1792_inR65;
  logic [127:0] zll_main_multiply1792_outR65;
  logic [256:0] zll_main_multiply1749_inR31;
  logic [127:0] zll_main_multiply1749_outR31;
  logic [383:0] zll_main_multiply300_in;
  logic [127:0] id_inR197;
  logic [0:0] rewire_prelude_not_inR65;
  logic [0:0] rewire_prelude_not_outR65;
  logic [128:0] zll_main_multiply1785_inR65;
  logic [127:0] zll_main_multiply1785_outR65;
  logic [383:0] zll_main_multiply1709_in;
  logic [127:0] id_inR198;
  logic [384:0] zll_main_multiply1_in;
  logic [127:0] id_inR199;
  logic [128:0] zll_main_multiply1792_inR66;
  logic [127:0] zll_main_multiply1792_outR66;
  logic [256:0] zll_main_multiply1788_inR34;
  logic [127:0] zll_main_multiply1788_outR34;
  logic [383:0] zll_main_multiply837_in;
  logic [127:0] id_inR200;
  logic [0:0] rewire_prelude_not_inR66;
  logic [0:0] rewire_prelude_not_outR66;
  logic [128:0] zll_main_multiply1785_inR66;
  logic [127:0] zll_main_multiply1785_outR66;
  logic [383:0] zll_main_multiply714_in;
  logic [127:0] id_inR201;
  logic [384:0] zll_main_multiply1098_in;
  logic [127:0] id_inR202;
  logic [128:0] zll_main_multiply1792_inR67;
  logic [127:0] zll_main_multiply1792_outR67;
  logic [256:0] zll_main_multiply1749_inR32;
  logic [127:0] zll_main_multiply1749_outR32;
  logic [383:0] zll_main_multiply940_in;
  logic [127:0] id_inR203;
  logic [0:0] rewire_prelude_not_inR67;
  logic [0:0] rewire_prelude_not_outR67;
  logic [128:0] zll_main_multiply1785_inR67;
  logic [127:0] zll_main_multiply1785_outR67;
  logic [383:0] zll_main_multiply76_in;
  logic [127:0] id_inR204;
  logic [384:0] zll_main_multiply344_in;
  logic [127:0] id_inR205;
  logic [128:0] zll_main_multiply1792_inR68;
  logic [127:0] zll_main_multiply1792_outR68;
  logic [256:0] zll_main_multiply1788_inR35;
  logic [127:0] zll_main_multiply1788_outR35;
  logic [383:0] zll_main_multiply970_in;
  logic [127:0] id_inR206;
  logic [0:0] rewire_prelude_not_inR68;
  logic [0:0] rewire_prelude_not_outR68;
  logic [128:0] zll_main_multiply1785_inR68;
  logic [127:0] zll_main_multiply1785_outR68;
  logic [383:0] zll_main_multiply1765_in;
  logic [127:0] id_inR207;
  logic [384:0] zll_main_multiply1336_in;
  logic [127:0] id_inR208;
  logic [128:0] zll_main_multiply1792_inR69;
  logic [127:0] zll_main_multiply1792_outR69;
  logic [256:0] zll_main_multiply1788_inR36;
  logic [127:0] zll_main_multiply1788_outR36;
  logic [383:0] zll_main_multiply1781_in;
  logic [127:0] id_inR209;
  logic [0:0] rewire_prelude_not_inR69;
  logic [0:0] rewire_prelude_not_outR69;
  logic [128:0] zll_main_multiply1785_inR69;
  logic [127:0] zll_main_multiply1785_outR69;
  logic [383:0] zll_main_multiply1657_in;
  logic [127:0] id_inR210;
  logic [384:0] zll_main_multiply630_in;
  logic [127:0] id_inR211;
  logic [128:0] zll_main_multiply1792_inR70;
  logic [127:0] zll_main_multiply1792_outR70;
  logic [256:0] zll_main_multiply1749_inR33;
  logic [127:0] zll_main_multiply1749_outR33;
  logic [383:0] zll_main_multiply1717_in;
  logic [127:0] id_inR212;
  logic [0:0] rewire_prelude_not_inR70;
  logic [0:0] rewire_prelude_not_outR70;
  logic [128:0] zll_main_multiply1785_inR70;
  logic [127:0] zll_main_multiply1785_outR70;
  logic [383:0] zll_main_multiply482_in;
  logic [127:0] id_inR213;
  logic [384:0] zll_main_multiply1158_in;
  logic [127:0] id_inR214;
  logic [128:0] zll_main_multiply1792_inR71;
  logic [127:0] zll_main_multiply1792_outR71;
  logic [256:0] zll_main_multiply1788_inR37;
  logic [127:0] zll_main_multiply1788_outR37;
  logic [383:0] zll_main_multiply281_in;
  logic [127:0] id_inR215;
  logic [0:0] rewire_prelude_not_inR71;
  logic [0:0] rewire_prelude_not_outR71;
  logic [128:0] zll_main_multiply1785_inR71;
  logic [127:0] zll_main_multiply1785_outR71;
  logic [383:0] zll_main_multiply1720_in;
  logic [127:0] id_inR216;
  logic [384:0] zll_main_multiply1640_in;
  logic [127:0] id_inR217;
  logic [128:0] zll_main_multiply1792_inR72;
  logic [127:0] zll_main_multiply1792_outR72;
  logic [256:0] zll_main_multiply1749_inR34;
  logic [127:0] zll_main_multiply1749_outR34;
  logic [383:0] zll_main_multiply268_in;
  logic [127:0] id_inR218;
  logic [0:0] rewire_prelude_not_inR72;
  logic [0:0] rewire_prelude_not_outR72;
  logic [128:0] zll_main_multiply1785_inR72;
  logic [127:0] zll_main_multiply1785_outR72;
  logic [383:0] zll_main_multiply603_in;
  logic [127:0] id_inR219;
  logic [384:0] zll_main_multiply55_in;
  logic [127:0] id_inR220;
  logic [128:0] zll_main_multiply1792_inR73;
  logic [127:0] zll_main_multiply1792_outR73;
  logic [256:0] zll_main_multiply1788_inR38;
  logic [127:0] zll_main_multiply1788_outR38;
  logic [383:0] zll_main_multiply23_in;
  logic [127:0] id_inR221;
  logic [0:0] rewire_prelude_not_inR73;
  logic [0:0] rewire_prelude_not_outR73;
  logic [128:0] zll_main_multiply1785_inR73;
  logic [127:0] zll_main_multiply1785_outR73;
  logic [383:0] zll_main_multiply1399_in;
  logic [127:0] id_inR222;
  logic [384:0] zll_main_multiply1637_in;
  logic [127:0] id_inR223;
  logic [128:0] zll_main_multiply1792_inR74;
  logic [127:0] zll_main_multiply1792_outR74;
  logic [256:0] zll_main_multiply1788_inR39;
  logic [127:0] zll_main_multiply1788_outR39;
  logic [383:0] zll_main_multiply1662_in;
  logic [127:0] id_inR224;
  logic [0:0] rewire_prelude_not_inR74;
  logic [0:0] rewire_prelude_not_outR74;
  logic [128:0] zll_main_multiply1785_inR74;
  logic [127:0] zll_main_multiply1785_outR74;
  logic [383:0] zll_main_multiply1106_in;
  logic [127:0] id_inR225;
  logic [384:0] zll_main_multiply1264_in;
  logic [127:0] id_inR226;
  logic [128:0] zll_main_multiply1792_inR75;
  logic [127:0] zll_main_multiply1792_outR75;
  logic [256:0] zll_main_multiply1788_inR40;
  logic [127:0] zll_main_multiply1788_outR40;
  logic [383:0] zll_main_multiply24_in;
  logic [127:0] id_inR227;
  logic [0:0] rewire_prelude_not_inR75;
  logic [0:0] rewire_prelude_not_outR75;
  logic [128:0] zll_main_multiply1785_inR75;
  logic [127:0] zll_main_multiply1785_outR75;
  logic [383:0] zll_main_multiply172_in;
  logic [127:0] id_inR228;
  logic [384:0] zll_main_multiply771_in;
  logic [127:0] id_inR229;
  logic [128:0] zll_main_multiply1792_inR76;
  logic [127:0] zll_main_multiply1792_outR76;
  logic [256:0] zll_main_multiply1788_inR41;
  logic [127:0] zll_main_multiply1788_outR41;
  logic [383:0] zll_main_multiply1587_in;
  logic [127:0] id_inR230;
  logic [0:0] rewire_prelude_not_inR76;
  logic [0:0] rewire_prelude_not_outR76;
  logic [128:0] zll_main_multiply1785_inR76;
  logic [127:0] zll_main_multiply1785_outR76;
  logic [383:0] zll_main_multiply1550_in;
  logic [127:0] id_inR231;
  logic [384:0] zll_main_multiply1167_in;
  logic [127:0] id_inR232;
  logic [128:0] zll_main_multiply1792_inR77;
  logic [127:0] zll_main_multiply1792_outR77;
  logic [256:0] zll_main_multiply1788_inR42;
  logic [127:0] zll_main_multiply1788_outR42;
  logic [383:0] zll_main_multiply1251_in;
  logic [127:0] id_inR233;
  logic [0:0] rewire_prelude_not_inR77;
  logic [0:0] rewire_prelude_not_outR77;
  logic [128:0] zll_main_multiply1785_inR77;
  logic [127:0] zll_main_multiply1785_outR77;
  logic [383:0] zll_main_multiply1320_in;
  logic [127:0] id_inR234;
  logic [384:0] zll_main_multiply43_in;
  logic [127:0] id_inR235;
  logic [128:0] zll_main_multiply1792_inR78;
  logic [127:0] zll_main_multiply1792_outR78;
  logic [256:0] zll_main_multiply1788_inR43;
  logic [127:0] zll_main_multiply1788_outR43;
  logic [383:0] zll_main_multiply1554_in;
  logic [127:0] id_inR236;
  logic [0:0] rewire_prelude_not_inR78;
  logic [0:0] rewire_prelude_not_outR78;
  logic [128:0] zll_main_multiply1785_inR78;
  logic [127:0] zll_main_multiply1785_outR78;
  logic [383:0] zll_main_multiply257_in;
  logic [127:0] id_inR237;
  logic [384:0] zll_main_multiply1513_in;
  logic [127:0] id_inR238;
  logic [128:0] zll_main_multiply1792_inR79;
  logic [127:0] zll_main_multiply1792_outR79;
  logic [256:0] zll_main_multiply1788_inR44;
  logic [127:0] zll_main_multiply1788_outR44;
  logic [383:0] zll_main_multiply113_in;
  logic [127:0] id_inR239;
  logic [0:0] rewire_prelude_not_inR79;
  logic [0:0] rewire_prelude_not_outR79;
  logic [128:0] zll_main_multiply1785_inR79;
  logic [127:0] zll_main_multiply1785_outR79;
  logic [383:0] zll_main_multiply1091_in;
  logic [127:0] id_inR240;
  logic [384:0] zll_main_multiply1266_in;
  logic [127:0] id_inR241;
  logic [128:0] zll_main_multiply1792_inR80;
  logic [127:0] zll_main_multiply1792_outR80;
  logic [256:0] zll_main_multiply1788_inR45;
  logic [127:0] zll_main_multiply1788_outR45;
  logic [383:0] zll_main_multiply418_in;
  logic [127:0] id_inR242;
  logic [0:0] rewire_prelude_not_inR80;
  logic [0:0] rewire_prelude_not_outR80;
  logic [128:0] zll_main_multiply1785_inR80;
  logic [127:0] zll_main_multiply1785_outR80;
  logic [383:0] zll_main_multiply409_in;
  logic [127:0] id_inR243;
  logic [384:0] zll_main_multiply726_in;
  logic [127:0] id_inR244;
  logic [128:0] zll_main_multiply1792_inR81;
  logic [127:0] zll_main_multiply1792_outR81;
  logic [256:0] zll_main_multiply1788_inR46;
  logic [127:0] zll_main_multiply1788_outR46;
  logic [383:0] zll_main_multiply1387_in;
  logic [127:0] id_inR245;
  logic [0:0] rewire_prelude_not_inR81;
  logic [0:0] rewire_prelude_not_outR81;
  logic [128:0] zll_main_multiply1785_inR81;
  logic [127:0] zll_main_multiply1785_outR81;
  logic [383:0] zll_main_multiply584_in;
  logic [127:0] id_inR246;
  logic [384:0] zll_main_multiply764_in;
  logic [127:0] id_inR247;
  logic [128:0] zll_main_multiply1792_inR82;
  logic [127:0] zll_main_multiply1792_outR82;
  logic [256:0] zll_main_multiply1788_inR47;
  logic [127:0] zll_main_multiply1788_outR47;
  logic [383:0] zll_main_multiply1627_in;
  logic [127:0] id_inR248;
  logic [0:0] rewire_prelude_not_inR82;
  logic [0:0] rewire_prelude_not_outR82;
  logic [128:0] zll_main_multiply1785_inR82;
  logic [127:0] zll_main_multiply1785_outR82;
  logic [383:0] zll_main_multiply442_in;
  logic [127:0] id_inR249;
  logic [384:0] zll_main_multiply1121_in;
  logic [127:0] id_inR250;
  logic [128:0] zll_main_multiply1792_inR83;
  logic [127:0] zll_main_multiply1792_outR83;
  logic [256:0] zll_main_multiply1788_inR48;
  logic [127:0] zll_main_multiply1788_outR48;
  logic [383:0] zll_main_multiply223_in;
  logic [127:0] id_inR251;
  logic [0:0] rewire_prelude_not_inR83;
  logic [0:0] rewire_prelude_not_outR83;
  logic [128:0] zll_main_multiply1785_inR83;
  logic [127:0] zll_main_multiply1785_outR83;
  logic [383:0] zll_main_multiply1410_in;
  logic [127:0] id_inR252;
  logic [384:0] zll_main_multiply1147_in;
  logic [127:0] id_inR253;
  logic [128:0] zll_main_multiply1792_inR84;
  logic [127:0] zll_main_multiply1792_outR84;
  logic [256:0] zll_main_multiply1788_inR49;
  logic [127:0] zll_main_multiply1788_outR49;
  logic [383:0] zll_main_multiply1137_in;
  logic [127:0] id_inR254;
  logic [0:0] rewire_prelude_not_inR84;
  logic [0:0] rewire_prelude_not_outR84;
  logic [128:0] zll_main_multiply1785_inR84;
  logic [127:0] zll_main_multiply1785_outR84;
  logic [383:0] zll_main_multiply1582_in;
  logic [127:0] id_inR255;
  logic [384:0] zll_main_multiply47_in;
  logic [127:0] id_inR256;
  logic [128:0] zll_main_multiply1792_inR85;
  logic [127:0] zll_main_multiply1792_outR85;
  logic [256:0] zll_main_multiply1749_inR35;
  logic [127:0] zll_main_multiply1749_outR35;
  logic [383:0] zll_main_multiply1047_in;
  logic [127:0] id_inR257;
  logic [0:0] rewire_prelude_not_inR85;
  logic [0:0] rewire_prelude_not_outR85;
  logic [128:0] zll_main_multiply1785_inR85;
  logic [127:0] zll_main_multiply1785_outR85;
  logic [383:0] zll_main_multiply98_in;
  logic [127:0] id_inR258;
  logic [384:0] zll_main_multiply1104_in;
  logic [127:0] id_inR259;
  logic [128:0] zll_main_multiply1792_inR86;
  logic [127:0] zll_main_multiply1792_outR86;
  logic [256:0] zll_main_multiply1749_inR36;
  logic [127:0] zll_main_multiply1749_outR36;
  logic [383:0] zll_main_multiply345_in;
  logic [127:0] id_inR260;
  logic [0:0] rewire_prelude_not_inR86;
  logic [0:0] rewire_prelude_not_outR86;
  logic [128:0] zll_main_multiply1785_inR86;
  logic [127:0] zll_main_multiply1785_outR86;
  logic [383:0] zll_main_multiply1438_in;
  logic [127:0] id_inR261;
  logic [384:0] zll_main_multiply1483_in;
  logic [127:0] id_inR262;
  logic [128:0] zll_main_multiply1792_inR87;
  logic [127:0] zll_main_multiply1792_outR87;
  logic [256:0] zll_main_multiply1788_inR50;
  logic [127:0] zll_main_multiply1788_outR50;
  logic [383:0] zll_main_multiply56_in;
  logic [127:0] id_inR263;
  logic [0:0] rewire_prelude_not_inR87;
  logic [0:0] rewire_prelude_not_outR87;
  logic [128:0] zll_main_multiply1785_inR87;
  logic [127:0] zll_main_multiply1785_outR87;
  logic [383:0] zll_main_multiply1200_in;
  logic [127:0] id_inR264;
  logic [384:0] zll_main_multiply800_in;
  logic [127:0] id_inR265;
  logic [128:0] zll_main_multiply1792_inR88;
  logic [127:0] zll_main_multiply1792_outR88;
  logic [256:0] zll_main_multiply1788_inR51;
  logic [127:0] zll_main_multiply1788_outR51;
  logic [383:0] zll_main_multiply411_in;
  logic [127:0] id_inR266;
  logic [0:0] rewire_prelude_not_inR88;
  logic [0:0] rewire_prelude_not_outR88;
  logic [128:0] zll_main_multiply1785_inR88;
  logic [127:0] zll_main_multiply1785_outR88;
  logic [383:0] zll_main_multiply774_in;
  logic [127:0] id_inR267;
  logic [384:0] zll_main_multiply129_in;
  logic [127:0] id_inR268;
  logic [128:0] zll_main_multiply1792_inR89;
  logic [127:0] zll_main_multiply1792_outR89;
  logic [256:0] zll_main_multiply1788_inR52;
  logic [127:0] zll_main_multiply1788_outR52;
  logic [383:0] zll_main_multiply1583_in;
  logic [127:0] id_inR269;
  logic [0:0] rewire_prelude_not_inR89;
  logic [0:0] rewire_prelude_not_outR89;
  logic [128:0] zll_main_multiply1785_inR89;
  logic [127:0] zll_main_multiply1785_outR89;
  logic [383:0] zll_main_multiply226_in;
  logic [127:0] id_inR270;
  logic [384:0] zll_main_multiply434_in;
  logic [127:0] id_inR271;
  logic [128:0] zll_main_multiply1792_inR90;
  logic [127:0] zll_main_multiply1792_outR90;
  logic [256:0] zll_main_multiply1788_inR53;
  logic [127:0] zll_main_multiply1788_outR53;
  logic [383:0] zll_main_multiply1369_in;
  logic [127:0] id_inR272;
  logic [0:0] rewire_prelude_not_inR90;
  logic [0:0] rewire_prelude_not_outR90;
  logic [128:0] zll_main_multiply1785_inR90;
  logic [127:0] zll_main_multiply1785_outR90;
  logic [383:0] zll_main_multiply697_in;
  logic [127:0] id_inR273;
  logic [384:0] zll_main_multiply869_in;
  logic [127:0] id_inR274;
  logic [128:0] zll_main_multiply1792_inR91;
  logic [127:0] zll_main_multiply1792_outR91;
  logic [256:0] zll_main_multiply1788_inR54;
  logic [127:0] zll_main_multiply1788_outR54;
  logic [383:0] zll_main_multiply1774_in;
  logic [127:0] id_inR275;
  logic [0:0] rewire_prelude_not_inR91;
  logic [0:0] rewire_prelude_not_outR91;
  logic [128:0] zll_main_multiply1785_inR91;
  logic [127:0] zll_main_multiply1785_outR91;
  logic [383:0] zll_main_multiply779_in;
  logic [127:0] id_inR276;
  logic [384:0] zll_main_multiply1551_in;
  logic [127:0] id_inR277;
  logic [128:0] zll_main_multiply1792_inR92;
  logic [127:0] zll_main_multiply1792_outR92;
  logic [256:0] zll_main_multiply1749_inR37;
  logic [127:0] zll_main_multiply1749_outR37;
  logic [383:0] zll_main_multiply845_in;
  logic [127:0] id_inR278;
  logic [0:0] rewire_prelude_not_inR92;
  logic [0:0] rewire_prelude_not_outR92;
  logic [128:0] zll_main_multiply1785_inR92;
  logic [127:0] zll_main_multiply1785_outR92;
  logic [383:0] zll_main_multiply565_in;
  logic [127:0] id_inR279;
  logic [384:0] zll_main_multiply496_in;
  logic [127:0] id_inR280;
  logic [128:0] zll_main_multiply1792_inR93;
  logic [127:0] zll_main_multiply1792_outR93;
  logic [256:0] zll_main_multiply1788_inR55;
  logic [127:0] zll_main_multiply1788_outR55;
  logic [383:0] zll_main_multiply1479_in;
  logic [127:0] id_inR281;
  logic [0:0] rewire_prelude_not_inR93;
  logic [0:0] rewire_prelude_not_outR93;
  logic [128:0] zll_main_multiply1785_inR93;
  logic [127:0] zll_main_multiply1785_outR93;
  logic [383:0] zll_main_multiply703_in;
  logic [127:0] id_inR282;
  logic [384:0] zll_main_multiply1286_in;
  logic [127:0] id_inR283;
  logic [128:0] zll_main_multiply1792_inR94;
  logic [127:0] zll_main_multiply1792_outR94;
  logic [256:0] zll_main_multiply1749_inR38;
  logic [127:0] zll_main_multiply1749_outR38;
  logic [383:0] zll_main_multiply293_in;
  logic [127:0] id_inR284;
  logic [0:0] rewire_prelude_not_inR94;
  logic [0:0] rewire_prelude_not_outR94;
  logic [128:0] zll_main_multiply1785_inR94;
  logic [127:0] zll_main_multiply1785_outR94;
  logic [383:0] zll_main_multiply1290_in;
  logic [127:0] id_inR285;
  logic [384:0] zll_main_multiply1189_in;
  logic [127:0] id_inR286;
  logic [128:0] zll_main_multiply1792_inR95;
  logic [127:0] zll_main_multiply1792_outR95;
  logic [256:0] zll_main_multiply1788_inR56;
  logic [127:0] zll_main_multiply1788_outR56;
  logic [383:0] zll_main_multiply1404_in;
  logic [127:0] id_inR287;
  logic [0:0] rewire_prelude_not_inR95;
  logic [0:0] rewire_prelude_not_outR95;
  logic [128:0] zll_main_multiply1785_inR95;
  logic [127:0] zll_main_multiply1785_outR95;
  logic [383:0] zll_main_multiply676_in;
  logic [127:0] id_inR288;
  logic [384:0] zll_main_multiply1769_in;
  logic [127:0] id_inR289;
  logic [128:0] zll_main_multiply1792_inR96;
  logic [127:0] zll_main_multiply1792_outR96;
  logic [256:0] zll_main_multiply1788_inR57;
  logic [127:0] zll_main_multiply1788_outR57;
  logic [383:0] zll_main_multiply464_in;
  logic [127:0] id_inR290;
  logic [0:0] rewire_prelude_not_inR96;
  logic [0:0] rewire_prelude_not_outR96;
  logic [128:0] zll_main_multiply1785_inR96;
  logic [127:0] zll_main_multiply1785_outR96;
  logic [383:0] zll_main_multiply538_in;
  logic [127:0] id_inR291;
  logic [384:0] zll_main_multiply175_in;
  logic [127:0] id_inR292;
  logic [128:0] zll_main_multiply1792_inR97;
  logic [127:0] zll_main_multiply1792_outR97;
  logic [256:0] zll_main_multiply1749_inR39;
  logic [127:0] zll_main_multiply1749_outR39;
  logic [383:0] zll_main_multiply376_in;
  logic [127:0] id_inR293;
  logic [0:0] rewire_prelude_not_inR97;
  logic [0:0] rewire_prelude_not_outR97;
  logic [128:0] zll_main_multiply1785_inR97;
  logic [127:0] zll_main_multiply1785_outR97;
  logic [383:0] zll_main_multiply471_in;
  logic [127:0] id_inR294;
  logic [384:0] zll_main_multiply872_in;
  logic [127:0] id_inR295;
  logic [128:0] zll_main_multiply1792_inR98;
  logic [127:0] zll_main_multiply1792_outR98;
  logic [256:0] zll_main_multiply1788_inR58;
  logic [127:0] zll_main_multiply1788_outR58;
  logic [383:0] zll_main_multiply1031_in;
  logic [127:0] id_inR296;
  logic [0:0] rewire_prelude_not_inR98;
  logic [0:0] rewire_prelude_not_outR98;
  logic [128:0] zll_main_multiply1785_inR98;
  logic [127:0] zll_main_multiply1785_outR98;
  logic [383:0] zll_main_multiply639_in;
  logic [127:0] id_inR297;
  logic [384:0] zll_main_multiply401_in;
  logic [127:0] id_inR298;
  logic [128:0] zll_main_multiply1792_inR99;
  logic [127:0] zll_main_multiply1792_outR99;
  logic [256:0] zll_main_multiply1749_inR40;
  logic [127:0] zll_main_multiply1749_outR40;
  logic [383:0] zll_main_multiply1588_in;
  logic [127:0] id_inR299;
  logic [0:0] rewire_prelude_not_inR99;
  logic [0:0] rewire_prelude_not_outR99;
  logic [128:0] zll_main_multiply1785_inR99;
  logic [127:0] zll_main_multiply1785_outR99;
  logic [383:0] zll_main_multiply1029_in;
  logic [127:0] id_inR300;
  logic [384:0] zll_main_multiply1340_in;
  logic [127:0] id_inR301;
  logic [128:0] zll_main_multiply1792_inR100;
  logic [127:0] zll_main_multiply1792_outR100;
  logic [256:0] zll_main_multiply1788_inR59;
  logic [127:0] zll_main_multiply1788_outR59;
  logic [383:0] zll_main_multiply1080_in;
  logic [127:0] id_inR302;
  logic [0:0] rewire_prelude_not_inR100;
  logic [0:0] rewire_prelude_not_outR100;
  logic [128:0] zll_main_multiply1785_inR100;
  logic [127:0] zll_main_multiply1785_outR100;
  logic [383:0] zll_main_multiply988_in;
  logic [127:0] id_inR303;
  logic [384:0] zll_main_multiply1510_in;
  logic [127:0] id_inR304;
  logic [128:0] zll_main_multiply1792_inR101;
  logic [127:0] zll_main_multiply1792_outR101;
  logic [256:0] zll_main_multiply1749_inR41;
  logic [127:0] zll_main_multiply1749_outR41;
  logic [383:0] zll_main_multiply137_in;
  logic [127:0] id_inR305;
  logic [0:0] rewire_prelude_not_inR101;
  logic [0:0] rewire_prelude_not_outR101;
  logic [128:0] zll_main_multiply1785_inR101;
  logic [127:0] zll_main_multiply1785_outR101;
  logic [383:0] zll_main_multiply67_in;
  logic [127:0] id_inR306;
  logic [384:0] zll_main_multiply1678_in;
  logic [127:0] id_inR307;
  logic [128:0] zll_main_multiply1792_inR102;
  logic [127:0] zll_main_multiply1792_outR102;
  logic [256:0] zll_main_multiply1788_inR60;
  logic [127:0] zll_main_multiply1788_outR60;
  logic [383:0] zll_main_multiply662_in;
  logic [127:0] id_inR308;
  logic [0:0] rewire_prelude_not_inR102;
  logic [0:0] rewire_prelude_not_outR102;
  logic [128:0] zll_main_multiply1785_inR102;
  logic [127:0] zll_main_multiply1785_outR102;
  logic [383:0] zll_main_multiply319_in;
  logic [127:0] id_inR309;
  logic [384:0] zll_main_multiply817_in;
  logic [127:0] id_inR310;
  logic [128:0] zll_main_multiply1792_inR103;
  logic [127:0] zll_main_multiply1792_outR103;
  logic [256:0] zll_main_multiply1749_inR42;
  logic [127:0] zll_main_multiply1749_outR42;
  logic [383:0] zll_main_multiply2_in;
  logic [127:0] id_inR311;
  logic [0:0] rewire_prelude_not_inR103;
  logic [0:0] rewire_prelude_not_outR103;
  logic [128:0] zll_main_multiply1785_inR103;
  logic [127:0] zll_main_multiply1785_outR103;
  logic [383:0] zll_main_multiply912_in;
  logic [127:0] id_inR312;
  logic [384:0] zll_main_multiply1624_in;
  logic [127:0] id_inR313;
  logic [128:0] zll_main_multiply1792_inR104;
  logic [127:0] zll_main_multiply1792_outR104;
  logic [256:0] zll_main_multiply1749_inR43;
  logic [127:0] zll_main_multiply1749_outR43;
  logic [383:0] zll_main_multiply977_in;
  logic [127:0] id_inR314;
  logic [0:0] rewire_prelude_not_inR104;
  logic [0:0] rewire_prelude_not_outR104;
  logic [128:0] zll_main_multiply1785_inR104;
  logic [127:0] zll_main_multiply1785_outR104;
  logic [383:0] zll_main_multiply180_in;
  logic [127:0] id_inR315;
  logic [384:0] zll_main_multiply476_in;
  logic [127:0] id_inR316;
  logic [128:0] zll_main_multiply1792_inR105;
  logic [127:0] zll_main_multiply1792_outR105;
  logic [256:0] zll_main_multiply1749_inR44;
  logic [127:0] zll_main_multiply1749_outR44;
  logic [383:0] zll_main_multiply1599_in;
  logic [127:0] id_inR317;
  logic [0:0] rewire_prelude_not_inR105;
  logic [0:0] rewire_prelude_not_outR105;
  logic [128:0] zll_main_multiply1785_inR105;
  logic [127:0] zll_main_multiply1785_outR105;
  logic [383:0] zll_main_multiply255_in;
  logic [127:0] id_inR318;
  logic [384:0] zll_main_multiply1531_in;
  logic [127:0] id_inR319;
  logic [128:0] zll_main_multiply1792_inR106;
  logic [127:0] zll_main_multiply1792_outR106;
  logic [256:0] zll_main_multiply1749_inR45;
  logic [127:0] zll_main_multiply1749_outR45;
  logic [383:0] zll_main_multiply1083_in;
  logic [127:0] id_inR320;
  logic [0:0] rewire_prelude_not_inR106;
  logic [0:0] rewire_prelude_not_outR106;
  logic [128:0] zll_main_multiply1785_inR106;
  logic [127:0] zll_main_multiply1785_outR106;
  logic [383:0] zll_main_multiply989_in;
  logic [127:0] id_inR321;
  logic [384:0] zll_main_multiply947_in;
  logic [127:0] id_inR322;
  logic [128:0] zll_main_multiply1792_inR107;
  logic [127:0] zll_main_multiply1792_outR107;
  logic [256:0] zll_main_multiply1749_inR46;
  logic [127:0] zll_main_multiply1749_outR46;
  logic [383:0] zll_main_multiply1245_in;
  logic [127:0] id_inR323;
  logic [0:0] rewire_prelude_not_inR107;
  logic [0:0] rewire_prelude_not_outR107;
  logic [128:0] zll_main_multiply1785_inR107;
  logic [127:0] zll_main_multiply1785_outR107;
  logic [383:0] zll_main_multiply167_in;
  logic [127:0] id_inR324;
  logic [384:0] zll_main_multiply1045_in;
  logic [127:0] id_inR325;
  logic [128:0] zll_main_multiply1792_inR108;
  logic [127:0] zll_main_multiply1792_outR108;
  logic [256:0] zll_main_multiply1749_inR47;
  logic [127:0] zll_main_multiply1749_outR47;
  logic [383:0] zll_main_multiply348_in;
  logic [127:0] id_inR326;
  logic [0:0] rewire_prelude_not_inR108;
  logic [0:0] rewire_prelude_not_outR108;
  logic [128:0] zll_main_multiply1785_inR108;
  logic [127:0] zll_main_multiply1785_outR108;
  logic [383:0] zll_main_multiply444_in;
  logic [127:0] id_inR327;
  logic [384:0] zll_main_multiply19_in;
  logic [127:0] id_inR328;
  logic [128:0] zll_main_multiply1792_inR109;
  logic [127:0] zll_main_multiply1792_outR109;
  logic [256:0] zll_main_multiply1788_inR61;
  logic [127:0] zll_main_multiply1788_outR61;
  logic [383:0] zll_main_multiply130_in;
  logic [127:0] id_inR329;
  logic [0:0] rewire_prelude_not_inR109;
  logic [0:0] rewire_prelude_not_outR109;
  logic [128:0] zll_main_multiply1785_inR109;
  logic [127:0] zll_main_multiply1785_outR109;
  logic [383:0] zll_main_multiply1403_in;
  logic [127:0] id_inR330;
  logic [384:0] zll_main_multiply1323_in;
  logic [127:0] id_inR331;
  logic [128:0] zll_main_multiply1792_inR110;
  logic [127:0] zll_main_multiply1792_outR110;
  logic [256:0] zll_main_multiply1749_inR48;
  logic [127:0] zll_main_multiply1749_outR48;
  logic [383:0] zll_main_multiply1329_in;
  logic [127:0] id_inR332;
  logic [0:0] rewire_prelude_not_inR110;
  logic [0:0] rewire_prelude_not_outR110;
  logic [128:0] zll_main_multiply1785_inR110;
  logic [127:0] zll_main_multiply1785_outR110;
  logic [383:0] zll_main_multiply389_in;
  logic [127:0] id_inR333;
  logic [384:0] zll_main_multiply294_in;
  logic [127:0] id_inR334;
  logic [128:0] zll_main_multiply1792_inR111;
  logic [127:0] zll_main_multiply1792_outR111;
  logic [256:0] zll_main_multiply1749_inR49;
  logic [127:0] zll_main_multiply1749_outR49;
  logic [383:0] zll_main_multiply335_in;
  logic [127:0] id_inR335;
  logic [0:0] rewire_prelude_not_inR111;
  logic [0:0] rewire_prelude_not_outR111;
  logic [128:0] zll_main_multiply1785_inR111;
  logic [127:0] zll_main_multiply1785_outR111;
  logic [383:0] zll_main_multiply295_in;
  logic [127:0] id_inR336;
  logic [384:0] zll_main_multiply563_in;
  logic [127:0] id_inR337;
  logic [128:0] zll_main_multiply1792_inR112;
  logic [127:0] zll_main_multiply1792_outR112;
  logic [256:0] zll_main_multiply1749_inR50;
  logic [127:0] zll_main_multiply1749_outR50;
  logic [383:0] zll_main_multiply1696_in;
  logic [127:0] id_inR338;
  logic [0:0] rewire_prelude_not_inR112;
  logic [0:0] rewire_prelude_not_outR112;
  logic [128:0] zll_main_multiply1785_inR112;
  logic [127:0] zll_main_multiply1785_outR112;
  logic [383:0] zll_main_multiply1154_in;
  logic [127:0] id_inR339;
  logic [384:0] zll_main_multiply1017_in;
  logic [127:0] id_inR340;
  logic [128:0] zll_main_multiply1792_inR113;
  logic [127:0] zll_main_multiply1792_outR113;
  logic [256:0] zll_main_multiply1788_inR62;
  logic [127:0] zll_main_multiply1788_outR62;
  logic [383:0] zll_main_multiply1568_in;
  logic [127:0] id_inR341;
  logic [0:0] rewire_prelude_not_inR113;
  logic [0:0] rewire_prelude_not_outR113;
  logic [128:0] zll_main_multiply1785_inR113;
  logic [127:0] zll_main_multiply1785_outR113;
  logic [383:0] zll_main_multiply921_in;
  logic [127:0] id_inR342;
  logic [384:0] zll_main_multiply576_in;
  logic [127:0] id_inR343;
  logic [128:0] zll_main_multiply1792_inR114;
  logic [127:0] zll_main_multiply1792_outR114;
  logic [256:0] zll_main_multiply1749_inR51;
  logic [127:0] zll_main_multiply1749_outR51;
  logic [383:0] zll_main_multiply1358_in;
  logic [127:0] id_inR344;
  logic [0:0] rewire_prelude_not_inR114;
  logic [0:0] rewire_prelude_not_outR114;
  logic [128:0] zll_main_multiply1785_inR114;
  logic [127:0] zll_main_multiply1785_outR114;
  logic [383:0] zll_main_multiply606_in;
  logic [127:0] id_inR345;
  logic [384:0] zll_main_multiply567_in;
  logic [127:0] id_inR346;
  logic [128:0] zll_main_multiply1792_inR115;
  logic [127:0] zll_main_multiply1792_outR115;
  logic [256:0] zll_main_multiply1749_inR52;
  logic [127:0] zll_main_multiply1749_outR52;
  logic [383:0] zll_main_multiply793_in;
  logic [127:0] id_inR347;
  logic [0:0] rewire_prelude_not_inR115;
  logic [0:0] rewire_prelude_not_outR115;
  logic [128:0] zll_main_multiply1785_inR115;
  logic [127:0] zll_main_multiply1785_outR115;
  logic [383:0] zll_main_multiply636_in;
  logic [127:0] id_inR348;
  logic [384:0] zll_main_multiply299_in;
  logic [127:0] id_inR349;
  logic [128:0] zll_main_multiply1792_inR116;
  logic [127:0] zll_main_multiply1792_outR116;
  logic [256:0] zll_main_multiply1788_inR63;
  logic [127:0] zll_main_multiply1788_outR63;
  logic [383:0] zll_main_multiply1705_in;
  logic [127:0] id_inR350;
  logic [0:0] rewire_prelude_not_inR116;
  logic [0:0] rewire_prelude_not_outR116;
  logic [128:0] zll_main_multiply1785_inR116;
  logic [127:0] zll_main_multiply1785_outR116;
  logic [383:0] zll_main_multiply439_in;
  logic [127:0] id_inR351;
  logic [384:0] zll_main_multiply263_in;
  logic [127:0] id_inR352;
  logic [128:0] zll_main_multiply1792_inR117;
  logic [127:0] zll_main_multiply1792_outR117;
  logic [256:0] zll_main_multiply1788_inR64;
  logic [127:0] zll_main_multiply1788_outR64;
  logic [383:0] zll_main_multiply1220_in;
  logic [127:0] id_inR353;
  logic [0:0] rewire_prelude_not_inR117;
  logic [0:0] rewire_prelude_not_outR117;
  logic [128:0] zll_main_multiply1785_inR117;
  logic [127:0] zll_main_multiply1785_outR117;
  logic [383:0] zll_main_multiply430_in;
  logic [127:0] id_inR354;
  logic [384:0] zll_main_multiply930_in;
  logic [127:0] id_inR355;
  logic [128:0] zll_main_multiply1792_inR118;
  logic [127:0] zll_main_multiply1792_outR118;
  logic [256:0] zll_main_multiply1749_inR53;
  logic [127:0] zll_main_multiply1749_outR53;
  logic [383:0] zll_main_multiply443_in;
  logic [127:0] id_inR356;
  logic [0:0] rewire_prelude_not_inR118;
  logic [0:0] rewire_prelude_not_outR118;
  logic [128:0] zll_main_multiply1785_inR118;
  logic [127:0] zll_main_multiply1785_outR118;
  logic [383:0] zll_main_multiply515_in;
  logic [127:0] id_inR357;
  logic [384:0] zll_main_multiply763_in;
  logic [127:0] id_inR358;
  logic [128:0] zll_main_multiply1792_inR119;
  logic [127:0] zll_main_multiply1792_outR119;
  logic [256:0] zll_main_multiply1749_inR54;
  logic [127:0] zll_main_multiply1749_outR54;
  logic [383:0] zll_main_multiply1725_in;
  logic [127:0] id_inR359;
  logic [0:0] rewire_prelude_not_inR119;
  logic [0:0] rewire_prelude_not_outR119;
  logic [128:0] zll_main_multiply1785_inR119;
  logic [127:0] zll_main_multiply1785_outR119;
  logic [383:0] zll_main_multiply1425_in;
  logic [127:0] id_inR360;
  logic [384:0] zll_main_multiply1784_in;
  logic [127:0] id_inR361;
  logic [128:0] zll_main_multiply1792_inR120;
  logic [127:0] zll_main_multiply1792_outR120;
  logic [256:0] zll_main_multiply1749_inR55;
  logic [127:0] zll_main_multiply1749_outR55;
  logic [383:0] zll_main_multiply1306_in;
  logic [127:0] id_inR362;
  logic [0:0] rewire_prelude_not_inR120;
  logic [0:0] rewire_prelude_not_outR120;
  logic [128:0] zll_main_multiply1785_inR120;
  logic [127:0] zll_main_multiply1785_outR120;
  logic [383:0] zll_main_multiply1407_in;
  logic [127:0] id_inR363;
  logic [384:0] zll_main_multiply692_in;
  logic [127:0] id_inR364;
  logic [128:0] zll_main_multiply1792_inR121;
  logic [127:0] zll_main_multiply1792_outR121;
  logic [256:0] zll_main_multiply1788_inR65;
  logic [127:0] zll_main_multiply1788_outR65;
  logic [383:0] zll_main_multiply850_in;
  logic [127:0] id_inR365;
  logic [0:0] rewire_prelude_not_inR121;
  logic [0:0] rewire_prelude_not_outR121;
  logic [128:0] zll_main_multiply1785_inR121;
  logic [127:0] zll_main_multiply1785_outR121;
  logic [383:0] zll_main_multiply392_in;
  logic [127:0] id_inR366;
  logic [384:0] zll_main_multiply887_in;
  logic [127:0] id_inR367;
  logic [128:0] zll_main_multiply1792_inR122;
  logic [127:0] zll_main_multiply1792_outR122;
  logic [256:0] zll_main_multiply1788_inR66;
  logic [127:0] zll_main_multiply1788_outR66;
  logic [383:0] zll_main_multiply1426_in;
  logic [127:0] id_inR368;
  logic [0:0] rewire_prelude_not_inR122;
  logic [0:0] rewire_prelude_not_outR122;
  logic [128:0] zll_main_multiply1785_inR122;
  logic [127:0] zll_main_multiply1785_outR122;
  logic [383:0] zll_main_multiply1704_in;
  logic [127:0] id_inR369;
  logic [384:0] zll_main_multiply758_in;
  logic [127:0] id_inR370;
  logic [128:0] zll_main_multiply1792_inR123;
  logic [127:0] zll_main_multiply1792_outR123;
  logic [256:0] zll_main_multiply1749_inR56;
  logic [127:0] zll_main_multiply1749_outR56;
  logic [383:0] zll_main_multiply537_in;
  logic [127:0] id_inR371;
  logic [0:0] rewire_prelude_not_inR123;
  logic [0:0] rewire_prelude_not_outR123;
  logic [128:0] zll_main_multiply1785_inR123;
  logic [127:0] zll_main_multiply1785_outR123;
  logic [383:0] zll_main_multiply446_in;
  logic [127:0] id_inR372;
  logic [384:0] zll_main_multiply1681_in;
  logic [127:0] id_inR373;
  logic [128:0] zll_main_multiply1792_inR124;
  logic [127:0] zll_main_multiply1792_outR124;
  logic [256:0] zll_main_multiply1788_inR67;
  logic [127:0] zll_main_multiply1788_outR67;
  logic [383:0] zll_main_multiply1125_in;
  logic [127:0] id_inR374;
  logic [0:0] rewire_prelude_not_inR124;
  logic [0:0] rewire_prelude_not_outR124;
  logic [128:0] zll_main_multiply1785_inR124;
  logic [127:0] zll_main_multiply1785_outR124;
  logic [383:0] zll_main_multiply1429_in;
  logic [127:0] id_inR375;
  logic [384:0] zll_main_multiply881_in;
  logic [127:0] id_inR376;
  logic [128:0] zll_main_multiply1792_inR125;
  logic [127:0] zll_main_multiply1792_outR125;
  logic [256:0] zll_main_multiply1749_inR57;
  logic [127:0] zll_main_multiply1749_outR57;
  logic [383:0] zll_main_multiply1113_in;
  logic [127:0] id_inR377;
  logic [0:0] rewire_prelude_not_inR125;
  logic [0:0] rewire_prelude_not_outR125;
  logic [128:0] zll_main_multiply1785_inR125;
  logic [127:0] zll_main_multiply1785_outR125;
  logic [383:0] zll_main_multiply1192_in;
  logic [127:0] id_inR378;
  logic [384:0] zll_main_multiply695_in;
  logic [127:0] id_inR379;
  logic [128:0] zll_main_multiply1792_inR126;
  logic [127:0] zll_main_multiply1792_outR126;
  logic [256:0] zll_main_multiply1788_inR68;
  logic [127:0] zll_main_multiply1788_outR68;
  logic [383:0] zll_main_multiply360_in;
  logic [127:0] id_inR380;
  logic [0:0] rewire_prelude_not_inR126;
  logic [0:0] rewire_prelude_not_outR126;
  logic [128:0] zll_main_multiply1785_inR126;
  logic [127:0] zll_main_multiply1785_outR126;
  logic [383:0] zll_main_multiply767_in;
  logic [127:0] id_inR381;
  logic [384:0] zll_main_multiply608_in;
  logic [127:0] id_inR382;
  logic [128:0] zll_main_multiply1792_inR127;
  logic [127:0] zll_main_multiply1792_outR127;
  logic [256:0] zll_main_multiply1788_inR69;
  logic [127:0] zll_main_multiply1788_outR69;
  logic [0:0] __continue;
  assign zll_main_multiplyfun1_in = {__in0, __in1};
  assign main_multiply_in = zll_main_multiplyfun1_in[255:0];
  assign zll_main_multiply1304_in = {main_multiply_in[255:128], main_multiply_in[127:0]};
  assign zll_main_multiply1066_in = zll_main_multiply1304_in[255:0];
  assign zll_main_multiply1727_in = {zll_main_multiply1066_in[127:0], zll_main_multiply1066_in[255:128]};
  assign zll_main_multiply459_in = {{8'h80{1'h0}}, zll_main_multiply1727_in[255:128], zll_main_multiply1727_in[127:0]};
  assign id_in = zll_main_multiply459_in[255:128];
  assign zll_main_multiply1476_in = {zll_main_multiply459_in[127:0], zll_main_multiply459_in[383:256], zll_main_multiply459_in[255:128], id_in[127]};
  assign id_inR1 = zll_main_multiply1476_in[128:1];
  assign zll_main_multiply1792_in = {zll_main_multiply1476_in[256:129], id_inR1[127]};
  ZLL_Main_multiply1792  inst (zll_main_multiply1792_in[128:1], zll_main_multiply1792_in[0], zll_main_multiply1792_out);
  assign zll_main_multiply1788_in = {zll_main_multiply1476_in[384:257], zll_main_multiply1476_in[256:129], zll_main_multiply1476_in[0]};
  ZLL_Main_multiply1788  instR1 (zll_main_multiply1788_in[256:129], zll_main_multiply1788_in[128:1], zll_main_multiply1788_out);
  assign zll_main_multiply939_in = {zll_main_multiply459_in[127:0], zll_main_multiply459_in[255:128], (zll_main_multiply1788_in[0] == 1'h1) ? zll_main_multiply1788_out : zll_main_multiply1792_out};
  assign id_inR2 = zll_main_multiply939_in[383:256];
  assign rewire_prelude_not_in = id_inR2[0];
  ReWire_Prelude_not  instR2 (rewire_prelude_not_in[0], rewire_prelude_not_out);
  assign zll_main_multiply1785_in = {zll_main_multiply939_in[383:256], rewire_prelude_not_out};
  ZLL_Main_multiply1785  instR3 (zll_main_multiply1785_in[128:1], zll_main_multiply1785_in[0], zll_main_multiply1785_out);
  assign zll_main_multiply62_in = {zll_main_multiply939_in[127:0], zll_main_multiply939_in[255:128], zll_main_multiply1785_out};
  assign id_inR3 = zll_main_multiply62_in[255:128];
  assign zll_main_multiply1570_in = {zll_main_multiply62_in[383:256], zll_main_multiply62_in[127:0], zll_main_multiply62_in[255:128], id_inR3[126]};
  assign id_inR4 = zll_main_multiply1570_in[128:1];
  assign zll_main_multiply1792_inR1 = {zll_main_multiply1570_in[384:257], id_inR4[126]};
  ZLL_Main_multiply1792  instR4 (zll_main_multiply1792_inR1[128:1], zll_main_multiply1792_inR1[0], zll_main_multiply1792_outR1);
  assign zll_main_multiply1749_in = {zll_main_multiply1570_in[384:257], zll_main_multiply1570_in[256:129], zll_main_multiply1570_in[0]};
  ZLL_Main_multiply1749  instR5 (zll_main_multiply1749_in[256:129], zll_main_multiply1749_in[128:1], zll_main_multiply1749_out);
  assign zll_main_multiply637_in = {zll_main_multiply62_in[127:0], zll_main_multiply62_in[255:128], (zll_main_multiply1749_in[0] == 1'h1) ? zll_main_multiply1749_out : zll_main_multiply1792_outR1};
  assign id_inR5 = zll_main_multiply637_in[383:256];
  assign rewire_prelude_not_inR1 = id_inR5[0];
  ReWire_Prelude_not  instR6 (rewire_prelude_not_inR1[0], rewire_prelude_not_outR1);
  assign zll_main_multiply1785_inR1 = {zll_main_multiply637_in[383:256], rewire_prelude_not_outR1};
  ZLL_Main_multiply1785  instR7 (zll_main_multiply1785_inR1[128:1], zll_main_multiply1785_inR1[0], zll_main_multiply1785_outR1);
  assign zll_main_multiply1342_in = {zll_main_multiply637_in[255:128], zll_main_multiply637_in[127:0], zll_main_multiply1785_outR1};
  assign id_inR6 = zll_main_multiply1342_in[383:256];
  assign zll_main_multiply811_in = {zll_main_multiply1342_in[127:0], zll_main_multiply1342_in[383:256], zll_main_multiply1342_in[255:128], id_inR6[125]};
  assign id_inR7 = zll_main_multiply811_in[256:129];
  assign zll_main_multiply1792_inR2 = {zll_main_multiply811_in[128:1], id_inR7[125]};
  ZLL_Main_multiply1792  instR8 (zll_main_multiply1792_inR2[128:1], zll_main_multiply1792_inR2[0], zll_main_multiply1792_outR2);
  assign zll_main_multiply1788_inR1 = {zll_main_multiply811_in[384:257], zll_main_multiply811_in[128:1], zll_main_multiply811_in[0]};
  ZLL_Main_multiply1788  instR9 (zll_main_multiply1788_inR1[256:129], zll_main_multiply1788_inR1[128:1], zll_main_multiply1788_outR1);
  assign zll_main_multiply681_in = {zll_main_multiply1342_in[127:0], zll_main_multiply1342_in[383:256], (zll_main_multiply1788_inR1[0] == 1'h1) ? zll_main_multiply1788_outR1 : zll_main_multiply1792_outR2};
  assign id_inR8 = zll_main_multiply681_in[383:256];
  assign rewire_prelude_not_inR2 = id_inR8[0];
  ReWire_Prelude_not  instR10 (rewire_prelude_not_inR2[0], rewire_prelude_not_outR2);
  assign zll_main_multiply1785_inR2 = {zll_main_multiply681_in[383:256], rewire_prelude_not_outR2};
  ZLL_Main_multiply1785  instR11 (zll_main_multiply1785_inR2[128:1], zll_main_multiply1785_inR2[0], zll_main_multiply1785_outR2);
  assign zll_main_multiply1772_in = {zll_main_multiply681_in[255:128], zll_main_multiply681_in[127:0], zll_main_multiply1785_outR2};
  assign id_inR9 = zll_main_multiply1772_in[383:256];
  assign zll_main_multiply322_in = {zll_main_multiply1772_in[383:256], zll_main_multiply1772_in[127:0], zll_main_multiply1772_in[255:128], id_inR9[124]};
  assign id_inR10 = zll_main_multiply322_in[384:257];
  assign zll_main_multiply1792_inR3 = {zll_main_multiply322_in[128:1], id_inR10[124]};
  ZLL_Main_multiply1792  instR12 (zll_main_multiply1792_inR3[128:1], zll_main_multiply1792_inR3[0], zll_main_multiply1792_outR3);
  assign zll_main_multiply1788_inR2 = {zll_main_multiply322_in[256:129], zll_main_multiply322_in[128:1], zll_main_multiply322_in[0]};
  ZLL_Main_multiply1788  instR13 (zll_main_multiply1788_inR2[256:129], zll_main_multiply1788_inR2[128:1], zll_main_multiply1788_outR2);
  assign zll_main_multiply864_in = {zll_main_multiply1772_in[383:256], zll_main_multiply1772_in[127:0], (zll_main_multiply1788_inR2[0] == 1'h1) ? zll_main_multiply1788_outR2 : zll_main_multiply1792_outR3};
  assign id_inR11 = zll_main_multiply864_in[255:128];
  assign rewire_prelude_not_inR3 = id_inR11[0];
  ReWire_Prelude_not  instR14 (rewire_prelude_not_inR3[0], rewire_prelude_not_outR3);
  assign zll_main_multiply1785_inR3 = {zll_main_multiply864_in[255:128], rewire_prelude_not_outR3};
  ZLL_Main_multiply1785  instR15 (zll_main_multiply1785_inR3[128:1], zll_main_multiply1785_inR3[0], zll_main_multiply1785_outR3);
  assign zll_main_multiply516_in = {zll_main_multiply864_in[383:256], zll_main_multiply864_in[127:0], zll_main_multiply1785_outR3};
  assign id_inR12 = zll_main_multiply516_in[383:256];
  assign zll_main_multiply1041_in = {zll_main_multiply516_in[383:256], zll_main_multiply516_in[255:128], zll_main_multiply516_in[127:0], id_inR12[123]};
  assign id_inR13 = zll_main_multiply1041_in[384:257];
  assign zll_main_multiply1792_inR4 = {zll_main_multiply1041_in[256:129], id_inR13[123]};
  ZLL_Main_multiply1792  instR16 (zll_main_multiply1792_inR4[128:1], zll_main_multiply1792_inR4[0], zll_main_multiply1792_outR4);
  assign zll_main_multiply1749_inR1 = {zll_main_multiply1041_in[256:129], zll_main_multiply1041_in[128:1], zll_main_multiply1041_in[0]};
  ZLL_Main_multiply1749  instR17 (zll_main_multiply1749_inR1[256:129], zll_main_multiply1749_inR1[128:1], zll_main_multiply1749_outR1);
  assign zll_main_multiply1038_in = {zll_main_multiply516_in[383:256], zll_main_multiply516_in[127:0], (zll_main_multiply1749_inR1[0] == 1'h1) ? zll_main_multiply1749_outR1 : zll_main_multiply1792_outR4};
  assign id_inR14 = zll_main_multiply1038_in[255:128];
  assign rewire_prelude_not_inR4 = id_inR14[0];
  ReWire_Prelude_not  instR18 (rewire_prelude_not_inR4[0], rewire_prelude_not_outR4);
  assign zll_main_multiply1785_inR4 = {zll_main_multiply1038_in[255:128], rewire_prelude_not_outR4};
  ZLL_Main_multiply1785  instR19 (zll_main_multiply1785_inR4[128:1], zll_main_multiply1785_inR4[0], zll_main_multiply1785_outR4);
  assign zll_main_multiply151_in = {zll_main_multiply1038_in[127:0], zll_main_multiply1038_in[383:256], zll_main_multiply1785_outR4};
  assign id_inR15 = zll_main_multiply151_in[255:128];
  assign zll_main_multiply909_in = {zll_main_multiply151_in[127:0], zll_main_multiply151_in[383:256], zll_main_multiply151_in[255:128], id_inR15[122]};
  assign id_inR16 = zll_main_multiply909_in[128:1];
  assign zll_main_multiply1792_inR5 = {zll_main_multiply909_in[256:129], id_inR16[122]};
  ZLL_Main_multiply1792  instR20 (zll_main_multiply1792_inR5[128:1], zll_main_multiply1792_inR5[0], zll_main_multiply1792_outR5);
  assign zll_main_multiply1788_inR3 = {zll_main_multiply909_in[384:257], zll_main_multiply909_in[256:129], zll_main_multiply909_in[0]};
  ZLL_Main_multiply1788  instR21 (zll_main_multiply1788_inR3[256:129], zll_main_multiply1788_inR3[128:1], zll_main_multiply1788_outR3);
  assign zll_main_multiply1491_in = {zll_main_multiply151_in[127:0], zll_main_multiply151_in[255:128], (zll_main_multiply1788_inR3[0] == 1'h1) ? zll_main_multiply1788_outR3 : zll_main_multiply1792_outR5};
  assign id_inR17 = zll_main_multiply1491_in[383:256];
  assign rewire_prelude_not_inR5 = id_inR17[0];
  ReWire_Prelude_not  instR22 (rewire_prelude_not_inR5[0], rewire_prelude_not_outR5);
  assign zll_main_multiply1785_inR5 = {zll_main_multiply1491_in[383:256], rewire_prelude_not_outR5};
  ZLL_Main_multiply1785  instR23 (zll_main_multiply1785_inR5[128:1], zll_main_multiply1785_inR5[0], zll_main_multiply1785_outR5);
  assign zll_main_multiply628_in = {zll_main_multiply1491_in[255:128], zll_main_multiply1491_in[127:0], zll_main_multiply1785_outR5};
  assign id_inR18 = zll_main_multiply628_in[383:256];
  assign zll_main_multiply1395_in = {zll_main_multiply628_in[127:0], zll_main_multiply628_in[383:256], zll_main_multiply628_in[255:128], id_inR18[121]};
  assign id_inR19 = zll_main_multiply1395_in[256:129];
  assign zll_main_multiply1792_inR6 = {zll_main_multiply1395_in[128:1], id_inR19[121]};
  ZLL_Main_multiply1792  instR24 (zll_main_multiply1792_inR6[128:1], zll_main_multiply1792_inR6[0], zll_main_multiply1792_outR6);
  assign zll_main_multiply1788_inR4 = {zll_main_multiply1395_in[384:257], zll_main_multiply1395_in[128:1], zll_main_multiply1395_in[0]};
  ZLL_Main_multiply1788  instR25 (zll_main_multiply1788_inR4[256:129], zll_main_multiply1788_inR4[128:1], zll_main_multiply1788_outR4);
  assign zll_main_multiply305_in = {zll_main_multiply628_in[127:0], zll_main_multiply628_in[383:256], (zll_main_multiply1788_inR4[0] == 1'h1) ? zll_main_multiply1788_outR4 : zll_main_multiply1792_outR6};
  assign id_inR20 = zll_main_multiply305_in[383:256];
  assign rewire_prelude_not_inR6 = id_inR20[0];
  ReWire_Prelude_not  instR26 (rewire_prelude_not_inR6[0], rewire_prelude_not_outR6);
  assign zll_main_multiply1785_inR6 = {zll_main_multiply305_in[383:256], rewire_prelude_not_outR6};
  ZLL_Main_multiply1785  instR27 (zll_main_multiply1785_inR6[128:1], zll_main_multiply1785_inR6[0], zll_main_multiply1785_outR6);
  assign zll_main_multiply667_in = {zll_main_multiply305_in[127:0], zll_main_multiply305_in[255:128], zll_main_multiply1785_outR6};
  assign id_inR21 = zll_main_multiply667_in[255:128];
  assign zll_main_multiply218_in = {zll_main_multiply667_in[383:256], zll_main_multiply667_in[255:128], zll_main_multiply667_in[127:0], id_inR21[120]};
  assign id_inR22 = zll_main_multiply218_in[256:129];
  assign zll_main_multiply1792_inR7 = {zll_main_multiply218_in[384:257], id_inR22[120]};
  ZLL_Main_multiply1792  instR28 (zll_main_multiply1792_inR7[128:1], zll_main_multiply1792_inR7[0], zll_main_multiply1792_outR7);
  assign zll_main_multiply1749_inR2 = {zll_main_multiply218_in[384:257], zll_main_multiply218_in[128:1], zll_main_multiply218_in[0]};
  ZLL_Main_multiply1749  instR29 (zll_main_multiply1749_inR2[256:129], zll_main_multiply1749_inR2[128:1], zll_main_multiply1749_outR2);
  assign zll_main_multiply97_in = {zll_main_multiply667_in[255:128], zll_main_multiply667_in[127:0], (zll_main_multiply1749_inR2[0] == 1'h1) ? zll_main_multiply1749_outR2 : zll_main_multiply1792_outR7};
  assign id_inR23 = zll_main_multiply97_in[255:128];
  assign rewire_prelude_not_inR7 = id_inR23[0];
  ReWire_Prelude_not  instR30 (rewire_prelude_not_inR7[0], rewire_prelude_not_outR7);
  assign zll_main_multiply1785_inR7 = {zll_main_multiply97_in[255:128], rewire_prelude_not_outR7};
  ZLL_Main_multiply1785  instR31 (zll_main_multiply1785_inR7[128:1], zll_main_multiply1785_inR7[0], zll_main_multiply1785_outR7);
  assign zll_main_multiply202_in = {zll_main_multiply97_in[127:0], zll_main_multiply97_in[383:256], zll_main_multiply1785_outR7};
  assign id_inR24 = zll_main_multiply202_in[255:128];
  assign zll_main_multiply143_in = {zll_main_multiply202_in[127:0], zll_main_multiply202_in[383:256], zll_main_multiply202_in[255:128], id_inR24[119]};
  assign id_inR25 = zll_main_multiply143_in[128:1];
  assign zll_main_multiply1792_inR8 = {zll_main_multiply143_in[256:129], id_inR25[119]};
  ZLL_Main_multiply1792  instR32 (zll_main_multiply1792_inR8[128:1], zll_main_multiply1792_inR8[0], zll_main_multiply1792_outR8);
  assign zll_main_multiply1788_inR5 = {zll_main_multiply143_in[384:257], zll_main_multiply143_in[256:129], zll_main_multiply143_in[0]};
  ZLL_Main_multiply1788  instR33 (zll_main_multiply1788_inR5[256:129], zll_main_multiply1788_inR5[128:1], zll_main_multiply1788_outR5);
  assign zll_main_multiply1630_in = {zll_main_multiply202_in[127:0], zll_main_multiply202_in[255:128], (zll_main_multiply1788_inR5[0] == 1'h1) ? zll_main_multiply1788_outR5 : zll_main_multiply1792_outR8};
  assign id_inR26 = zll_main_multiply1630_in[383:256];
  assign rewire_prelude_not_inR8 = id_inR26[0];
  ReWire_Prelude_not  instR34 (rewire_prelude_not_inR8[0], rewire_prelude_not_outR8);
  assign zll_main_multiply1785_inR8 = {zll_main_multiply1630_in[383:256], rewire_prelude_not_outR8};
  ZLL_Main_multiply1785  instR35 (zll_main_multiply1785_inR8[128:1], zll_main_multiply1785_inR8[0], zll_main_multiply1785_outR8);
  assign zll_main_multiply1766_in = {zll_main_multiply1630_in[127:0], zll_main_multiply1630_in[255:128], zll_main_multiply1785_outR8};
  assign id_inR27 = zll_main_multiply1766_in[255:128];
  assign zll_main_multiply918_in = {zll_main_multiply1766_in[127:0], zll_main_multiply1766_in[383:256], zll_main_multiply1766_in[255:128], id_inR27[118]};
  assign id_inR28 = zll_main_multiply918_in[128:1];
  assign zll_main_multiply1792_inR9 = {zll_main_multiply918_in[256:129], id_inR28[118]};
  ZLL_Main_multiply1792  instR36 (zll_main_multiply1792_inR9[128:1], zll_main_multiply1792_inR9[0], zll_main_multiply1792_outR9);
  assign zll_main_multiply1788_inR6 = {zll_main_multiply918_in[384:257], zll_main_multiply918_in[256:129], zll_main_multiply918_in[0]};
  ZLL_Main_multiply1788  instR37 (zll_main_multiply1788_inR6[256:129], zll_main_multiply1788_inR6[128:1], zll_main_multiply1788_outR6);
  assign zll_main_multiply978_in = {zll_main_multiply1766_in[127:0], zll_main_multiply1766_in[255:128], (zll_main_multiply1788_inR6[0] == 1'h1) ? zll_main_multiply1788_outR6 : zll_main_multiply1792_outR9};
  assign id_inR29 = zll_main_multiply978_in[383:256];
  assign rewire_prelude_not_inR9 = id_inR29[0];
  ReWire_Prelude_not  instR38 (rewire_prelude_not_inR9[0], rewire_prelude_not_outR9);
  assign zll_main_multiply1785_inR9 = {zll_main_multiply978_in[383:256], rewire_prelude_not_outR9};
  ZLL_Main_multiply1785  instR39 (zll_main_multiply1785_inR9[128:1], zll_main_multiply1785_inR9[0], zll_main_multiply1785_outR9);
  assign zll_main_multiply497_in = {zll_main_multiply978_in[127:0], zll_main_multiply978_in[255:128], zll_main_multiply1785_outR9};
  assign id_inR30 = zll_main_multiply497_in[255:128];
  assign zll_main_multiply617_in = {zll_main_multiply497_in[383:256], zll_main_multiply497_in[255:128], zll_main_multiply497_in[127:0], id_inR30[117]};
  assign id_inR31 = zll_main_multiply617_in[256:129];
  assign zll_main_multiply1792_inR10 = {zll_main_multiply617_in[384:257], id_inR31[117]};
  ZLL_Main_multiply1792  instR40 (zll_main_multiply1792_inR10[128:1], zll_main_multiply1792_inR10[0], zll_main_multiply1792_outR10);
  assign zll_main_multiply1749_inR3 = {zll_main_multiply617_in[384:257], zll_main_multiply617_in[128:1], zll_main_multiply617_in[0]};
  ZLL_Main_multiply1749  instR41 (zll_main_multiply1749_inR3[256:129], zll_main_multiply1749_inR3[128:1], zll_main_multiply1749_outR3);
  assign zll_main_multiply1473_in = {zll_main_multiply497_in[255:128], zll_main_multiply497_in[127:0], (zll_main_multiply1749_inR3[0] == 1'h1) ? zll_main_multiply1749_outR3 : zll_main_multiply1792_outR10};
  assign id_inR32 = zll_main_multiply1473_in[255:128];
  assign rewire_prelude_not_inR10 = id_inR32[0];
  ReWire_Prelude_not  instR42 (rewire_prelude_not_inR10[0], rewire_prelude_not_outR10);
  assign zll_main_multiply1785_inR10 = {zll_main_multiply1473_in[255:128], rewire_prelude_not_outR10};
  ZLL_Main_multiply1785  instR43 (zll_main_multiply1785_inR10[128:1], zll_main_multiply1785_inR10[0], zll_main_multiply1785_outR10);
  assign zll_main_multiply1206_in = {zll_main_multiply1473_in[383:256], zll_main_multiply1473_in[127:0], zll_main_multiply1785_outR10};
  assign id_inR33 = zll_main_multiply1206_in[383:256];
  assign zll_main_multiply158_in = {zll_main_multiply1206_in[383:256], zll_main_multiply1206_in[255:128], zll_main_multiply1206_in[127:0], id_inR33[116]};
  assign id_inR34 = zll_main_multiply158_in[384:257];
  assign zll_main_multiply1792_inR11 = {zll_main_multiply158_in[256:129], id_inR34[116]};
  ZLL_Main_multiply1792  instR44 (zll_main_multiply1792_inR11[128:1], zll_main_multiply1792_inR11[0], zll_main_multiply1792_outR11);
  assign zll_main_multiply1749_inR4 = {zll_main_multiply158_in[256:129], zll_main_multiply158_in[128:1], zll_main_multiply158_in[0]};
  ZLL_Main_multiply1749  instR45 (zll_main_multiply1749_inR4[256:129], zll_main_multiply1749_inR4[128:1], zll_main_multiply1749_outR4);
  assign zll_main_multiply769_in = {zll_main_multiply1206_in[383:256], zll_main_multiply1206_in[127:0], (zll_main_multiply1749_inR4[0] == 1'h1) ? zll_main_multiply1749_outR4 : zll_main_multiply1792_outR11};
  assign id_inR35 = zll_main_multiply769_in[255:128];
  assign rewire_prelude_not_inR11 = id_inR35[0];
  ReWire_Prelude_not  instR46 (rewire_prelude_not_inR11[0], rewire_prelude_not_outR11);
  assign zll_main_multiply1785_inR11 = {zll_main_multiply769_in[255:128], rewire_prelude_not_outR11};
  ZLL_Main_multiply1785  instR47 (zll_main_multiply1785_inR11[128:1], zll_main_multiply1785_inR11[0], zll_main_multiply1785_outR11);
  assign zll_main_multiply730_in = {zll_main_multiply769_in[127:0], zll_main_multiply769_in[383:256], zll_main_multiply1785_outR11};
  assign id_inR36 = zll_main_multiply730_in[255:128];
  assign zll_main_multiply1089_in = {zll_main_multiply730_in[383:256], zll_main_multiply730_in[127:0], zll_main_multiply730_in[255:128], id_inR36[115]};
  assign id_inR37 = zll_main_multiply1089_in[128:1];
  assign zll_main_multiply1792_inR12 = {zll_main_multiply1089_in[384:257], id_inR37[115]};
  ZLL_Main_multiply1792  instR48 (zll_main_multiply1792_inR12[128:1], zll_main_multiply1792_inR12[0], zll_main_multiply1792_outR12);
  assign zll_main_multiply1749_inR5 = {zll_main_multiply1089_in[384:257], zll_main_multiply1089_in[256:129], zll_main_multiply1089_in[0]};
  ZLL_Main_multiply1749  instR49 (zll_main_multiply1749_inR5[256:129], zll_main_multiply1749_inR5[128:1], zll_main_multiply1749_outR5);
  assign zll_main_multiply871_in = {zll_main_multiply730_in[127:0], zll_main_multiply730_in[255:128], (zll_main_multiply1749_inR5[0] == 1'h1) ? zll_main_multiply1749_outR5 : zll_main_multiply1792_outR12};
  assign id_inR38 = zll_main_multiply871_in[383:256];
  assign rewire_prelude_not_inR12 = id_inR38[0];
  ReWire_Prelude_not  instR50 (rewire_prelude_not_inR12[0], rewire_prelude_not_outR12);
  assign zll_main_multiply1785_inR12 = {zll_main_multiply871_in[383:256], rewire_prelude_not_outR12};
  ZLL_Main_multiply1785  instR51 (zll_main_multiply1785_inR12[128:1], zll_main_multiply1785_inR12[0], zll_main_multiply1785_outR12);
  assign zll_main_multiply279_in = {zll_main_multiply871_in[127:0], zll_main_multiply871_in[255:128], zll_main_multiply1785_outR12};
  assign id_inR39 = zll_main_multiply279_in[255:128];
  assign zll_main_multiply39_in = {zll_main_multiply279_in[383:256], zll_main_multiply279_in[127:0], zll_main_multiply279_in[255:128], id_inR39[114]};
  assign id_inR40 = zll_main_multiply39_in[128:1];
  assign zll_main_multiply1792_inR13 = {zll_main_multiply39_in[384:257], id_inR40[114]};
  ZLL_Main_multiply1792  instR52 (zll_main_multiply1792_inR13[128:1], zll_main_multiply1792_inR13[0], zll_main_multiply1792_outR13);
  assign zll_main_multiply1749_inR6 = {zll_main_multiply39_in[384:257], zll_main_multiply39_in[256:129], zll_main_multiply39_in[0]};
  ZLL_Main_multiply1749  instR53 (zll_main_multiply1749_inR6[256:129], zll_main_multiply1749_inR6[128:1], zll_main_multiply1749_outR6);
  assign zll_main_multiply1691_in = {zll_main_multiply279_in[127:0], zll_main_multiply279_in[255:128], (zll_main_multiply1749_inR6[0] == 1'h1) ? zll_main_multiply1749_outR6 : zll_main_multiply1792_outR13};
  assign id_inR41 = zll_main_multiply1691_in[383:256];
  assign rewire_prelude_not_inR13 = id_inR41[0];
  ReWire_Prelude_not  instR54 (rewire_prelude_not_inR13[0], rewire_prelude_not_outR13);
  assign zll_main_multiply1785_inR13 = {zll_main_multiply1691_in[383:256], rewire_prelude_not_outR13};
  ZLL_Main_multiply1785  instR55 (zll_main_multiply1785_inR13[128:1], zll_main_multiply1785_inR13[0], zll_main_multiply1785_outR13);
  assign zll_main_multiply1282_in = {zll_main_multiply1691_in[255:128], zll_main_multiply1691_in[127:0], zll_main_multiply1785_outR13};
  assign id_inR42 = zll_main_multiply1282_in[383:256];
  assign zll_main_multiply110_in = {zll_main_multiply1282_in[383:256], zll_main_multiply1282_in[255:128], zll_main_multiply1282_in[127:0], id_inR42[113]};
  assign id_inR43 = zll_main_multiply110_in[384:257];
  assign zll_main_multiply1792_inR14 = {zll_main_multiply110_in[256:129], id_inR43[113]};
  ZLL_Main_multiply1792  instR56 (zll_main_multiply1792_inR14[128:1], zll_main_multiply1792_inR14[0], zll_main_multiply1792_outR14);
  assign zll_main_multiply1749_inR7 = {zll_main_multiply110_in[256:129], zll_main_multiply110_in[128:1], zll_main_multiply110_in[0]};
  ZLL_Main_multiply1749  instR57 (zll_main_multiply1749_inR7[256:129], zll_main_multiply1749_inR7[128:1], zll_main_multiply1749_outR7);
  assign zll_main_multiply282_in = {zll_main_multiply1282_in[383:256], zll_main_multiply1282_in[127:0], (zll_main_multiply1749_inR7[0] == 1'h1) ? zll_main_multiply1749_outR7 : zll_main_multiply1792_outR14};
  assign id_inR44 = zll_main_multiply282_in[255:128];
  assign rewire_prelude_not_inR14 = id_inR44[0];
  ReWire_Prelude_not  instR58 (rewire_prelude_not_inR14[0], rewire_prelude_not_outR14);
  assign zll_main_multiply1785_inR14 = {zll_main_multiply282_in[255:128], rewire_prelude_not_outR14};
  ZLL_Main_multiply1785  instR59 (zll_main_multiply1785_inR14[128:1], zll_main_multiply1785_inR14[0], zll_main_multiply1785_outR14);
  assign zll_main_multiply71_in = {zll_main_multiply282_in[127:0], zll_main_multiply282_in[383:256], zll_main_multiply1785_outR14};
  assign id_inR45 = zll_main_multiply71_in[255:128];
  assign zll_main_multiply1176_in = {zll_main_multiply71_in[127:0], zll_main_multiply71_in[383:256], zll_main_multiply71_in[255:128], id_inR45[112]};
  assign id_inR46 = zll_main_multiply1176_in[128:1];
  assign zll_main_multiply1792_inR15 = {zll_main_multiply1176_in[256:129], id_inR46[112]};
  ZLL_Main_multiply1792  instR60 (zll_main_multiply1792_inR15[128:1], zll_main_multiply1792_inR15[0], zll_main_multiply1792_outR15);
  assign zll_main_multiply1788_inR7 = {zll_main_multiply1176_in[384:257], zll_main_multiply1176_in[256:129], zll_main_multiply1176_in[0]};
  ZLL_Main_multiply1788  instR61 (zll_main_multiply1788_inR7[256:129], zll_main_multiply1788_inR7[128:1], zll_main_multiply1788_outR7);
  assign zll_main_multiply910_in = {zll_main_multiply71_in[127:0], zll_main_multiply71_in[255:128], (zll_main_multiply1788_inR7[0] == 1'h1) ? zll_main_multiply1788_outR7 : zll_main_multiply1792_outR15};
  assign id_inR47 = zll_main_multiply910_in[383:256];
  assign rewire_prelude_not_inR15 = id_inR47[0];
  ReWire_Prelude_not  instR62 (rewire_prelude_not_inR15[0], rewire_prelude_not_outR15);
  assign zll_main_multiply1785_inR15 = {zll_main_multiply910_in[383:256], rewire_prelude_not_outR15};
  ZLL_Main_multiply1785  instR63 (zll_main_multiply1785_inR15[128:1], zll_main_multiply1785_inR15[0], zll_main_multiply1785_outR15);
  assign zll_main_multiply1165_in = {zll_main_multiply910_in[127:0], zll_main_multiply910_in[255:128], zll_main_multiply1785_outR15};
  assign id_inR48 = zll_main_multiply1165_in[255:128];
  assign zll_main_multiply168_in = {zll_main_multiply1165_in[127:0], zll_main_multiply1165_in[383:256], zll_main_multiply1165_in[255:128], id_inR48[111]};
  assign id_inR49 = zll_main_multiply168_in[128:1];
  assign zll_main_multiply1792_inR16 = {zll_main_multiply168_in[256:129], id_inR49[111]};
  ZLL_Main_multiply1792  instR64 (zll_main_multiply1792_inR16[128:1], zll_main_multiply1792_inR16[0], zll_main_multiply1792_outR16);
  assign zll_main_multiply1788_inR8 = {zll_main_multiply168_in[384:257], zll_main_multiply168_in[256:129], zll_main_multiply168_in[0]};
  ZLL_Main_multiply1788  instR65 (zll_main_multiply1788_inR8[256:129], zll_main_multiply1788_inR8[128:1], zll_main_multiply1788_outR8);
  assign zll_main_multiply195_in = {zll_main_multiply1165_in[127:0], zll_main_multiply1165_in[255:128], (zll_main_multiply1788_inR8[0] == 1'h1) ? zll_main_multiply1788_outR8 : zll_main_multiply1792_outR16};
  assign id_inR50 = zll_main_multiply195_in[383:256];
  assign rewire_prelude_not_inR16 = id_inR50[0];
  ReWire_Prelude_not  instR66 (rewire_prelude_not_inR16[0], rewire_prelude_not_outR16);
  assign zll_main_multiply1785_inR16 = {zll_main_multiply195_in[383:256], rewire_prelude_not_outR16};
  ZLL_Main_multiply1785  instR67 (zll_main_multiply1785_inR16[128:1], zll_main_multiply1785_inR16[0], zll_main_multiply1785_outR16);
  assign zll_main_multiply750_in = {zll_main_multiply195_in[127:0], zll_main_multiply195_in[255:128], zll_main_multiply1785_outR16};
  assign id_inR51 = zll_main_multiply750_in[255:128];
  assign zll_main_multiply196_in = {zll_main_multiply750_in[127:0], zll_main_multiply750_in[383:256], zll_main_multiply750_in[255:128], id_inR51[110]};
  assign id_inR52 = zll_main_multiply196_in[128:1];
  assign zll_main_multiply1792_inR17 = {zll_main_multiply196_in[256:129], id_inR52[110]};
  ZLL_Main_multiply1792  instR68 (zll_main_multiply1792_inR17[128:1], zll_main_multiply1792_inR17[0], zll_main_multiply1792_outR17);
  assign zll_main_multiply1788_inR9 = {zll_main_multiply196_in[384:257], zll_main_multiply196_in[256:129], zll_main_multiply196_in[0]};
  ZLL_Main_multiply1788  instR69 (zll_main_multiply1788_inR9[256:129], zll_main_multiply1788_inR9[128:1], zll_main_multiply1788_outR9);
  assign zll_main_multiply765_in = {zll_main_multiply750_in[127:0], zll_main_multiply750_in[255:128], (zll_main_multiply1788_inR9[0] == 1'h1) ? zll_main_multiply1788_outR9 : zll_main_multiply1792_outR17};
  assign id_inR53 = zll_main_multiply765_in[383:256];
  assign rewire_prelude_not_inR17 = id_inR53[0];
  ReWire_Prelude_not  instR70 (rewire_prelude_not_inR17[0], rewire_prelude_not_outR17);
  assign zll_main_multiply1785_inR17 = {zll_main_multiply765_in[383:256], rewire_prelude_not_outR17};
  ZLL_Main_multiply1785  instR71 (zll_main_multiply1785_inR17[128:1], zll_main_multiply1785_inR17[0], zll_main_multiply1785_outR17);
  assign zll_main_multiply851_in = {zll_main_multiply765_in[127:0], zll_main_multiply765_in[255:128], zll_main_multiply1785_outR17};
  assign id_inR54 = zll_main_multiply851_in[255:128];
  assign zll_main_multiply831_in = {zll_main_multiply851_in[127:0], zll_main_multiply851_in[383:256], zll_main_multiply851_in[255:128], id_inR54[109]};
  assign id_inR55 = zll_main_multiply831_in[128:1];
  assign zll_main_multiply1792_inR18 = {zll_main_multiply831_in[256:129], id_inR55[109]};
  ZLL_Main_multiply1792  instR72 (zll_main_multiply1792_inR18[128:1], zll_main_multiply1792_inR18[0], zll_main_multiply1792_outR18);
  assign zll_main_multiply1788_inR10 = {zll_main_multiply831_in[384:257], zll_main_multiply831_in[256:129], zll_main_multiply831_in[0]};
  ZLL_Main_multiply1788  instR73 (zll_main_multiply1788_inR10[256:129], zll_main_multiply1788_inR10[128:1], zll_main_multiply1788_outR10);
  assign zll_main_multiply1107_in = {zll_main_multiply851_in[127:0], zll_main_multiply851_in[255:128], (zll_main_multiply1788_inR10[0] == 1'h1) ? zll_main_multiply1788_outR10 : zll_main_multiply1792_outR18};
  assign id_inR56 = zll_main_multiply1107_in[383:256];
  assign rewire_prelude_not_inR18 = id_inR56[0];
  ReWire_Prelude_not  instR74 (rewire_prelude_not_inR18[0], rewire_prelude_not_outR18);
  assign zll_main_multiply1785_inR18 = {zll_main_multiply1107_in[383:256], rewire_prelude_not_outR18};
  ZLL_Main_multiply1785  instR75 (zll_main_multiply1785_inR18[128:1], zll_main_multiply1785_inR18[0], zll_main_multiply1785_outR18);
  assign zll_main_multiply29_in = {zll_main_multiply1107_in[255:128], zll_main_multiply1107_in[127:0], zll_main_multiply1785_outR18};
  assign id_inR57 = zll_main_multiply29_in[383:256];
  assign zll_main_multiply964_in = {zll_main_multiply29_in[127:0], zll_main_multiply29_in[383:256], zll_main_multiply29_in[255:128], id_inR57[108]};
  assign id_inR58 = zll_main_multiply964_in[256:129];
  assign zll_main_multiply1792_inR19 = {zll_main_multiply964_in[128:1], id_inR58[108]};
  ZLL_Main_multiply1792  instR76 (zll_main_multiply1792_inR19[128:1], zll_main_multiply1792_inR19[0], zll_main_multiply1792_outR19);
  assign zll_main_multiply1788_inR11 = {zll_main_multiply964_in[384:257], zll_main_multiply964_in[128:1], zll_main_multiply964_in[0]};
  ZLL_Main_multiply1788  instR77 (zll_main_multiply1788_inR11[256:129], zll_main_multiply1788_inR11[128:1], zll_main_multiply1788_outR11);
  assign zll_main_multiply1345_in = {zll_main_multiply29_in[127:0], zll_main_multiply29_in[383:256], (zll_main_multiply1788_inR11[0] == 1'h1) ? zll_main_multiply1788_outR11 : zll_main_multiply1792_outR19};
  assign id_inR59 = zll_main_multiply1345_in[383:256];
  assign rewire_prelude_not_inR19 = id_inR59[0];
  ReWire_Prelude_not  instR78 (rewire_prelude_not_inR19[0], rewire_prelude_not_outR19);
  assign zll_main_multiply1785_inR19 = {zll_main_multiply1345_in[383:256], rewire_prelude_not_outR19};
  ZLL_Main_multiply1785  instR79 (zll_main_multiply1785_inR19[128:1], zll_main_multiply1785_inR19[0], zll_main_multiply1785_outR19);
  assign zll_main_multiply390_in = {zll_main_multiply1345_in[255:128], zll_main_multiply1345_in[127:0], zll_main_multiply1785_outR19};
  assign id_inR60 = zll_main_multiply390_in[383:256];
  assign zll_main_multiply1076_in = {zll_main_multiply390_in[383:256], zll_main_multiply390_in[255:128], zll_main_multiply390_in[127:0], id_inR60[107]};
  assign id_inR61 = zll_main_multiply1076_in[384:257];
  assign zll_main_multiply1792_inR20 = {zll_main_multiply1076_in[256:129], id_inR61[107]};
  ZLL_Main_multiply1792  instR80 (zll_main_multiply1792_inR20[128:1], zll_main_multiply1792_inR20[0], zll_main_multiply1792_outR20);
  assign zll_main_multiply1749_inR8 = {zll_main_multiply1076_in[256:129], zll_main_multiply1076_in[128:1], zll_main_multiply1076_in[0]};
  ZLL_Main_multiply1749  instR81 (zll_main_multiply1749_inR8[256:129], zll_main_multiply1749_inR8[128:1], zll_main_multiply1749_outR8);
  assign zll_main_multiply687_in = {zll_main_multiply390_in[383:256], zll_main_multiply390_in[127:0], (zll_main_multiply1749_inR8[0] == 1'h1) ? zll_main_multiply1749_outR8 : zll_main_multiply1792_outR20};
  assign id_inR62 = zll_main_multiply687_in[255:128];
  assign rewire_prelude_not_inR20 = id_inR62[0];
  ReWire_Prelude_not  instR82 (rewire_prelude_not_inR20[0], rewire_prelude_not_outR20);
  assign zll_main_multiply1785_inR20 = {zll_main_multiply687_in[255:128], rewire_prelude_not_outR20};
  ZLL_Main_multiply1785  instR83 (zll_main_multiply1785_inR20[128:1], zll_main_multiply1785_inR20[0], zll_main_multiply1785_outR20);
  assign zll_main_multiply138_in = {zll_main_multiply687_in[383:256], zll_main_multiply687_in[127:0], zll_main_multiply1785_outR20};
  assign id_inR63 = zll_main_multiply138_in[383:256];
  assign zll_main_multiply1411_in = {zll_main_multiply138_in[383:256], zll_main_multiply138_in[127:0], zll_main_multiply138_in[255:128], id_inR63[106]};
  assign id_inR64 = zll_main_multiply1411_in[384:257];
  assign zll_main_multiply1792_inR21 = {zll_main_multiply1411_in[128:1], id_inR64[106]};
  ZLL_Main_multiply1792  instR84 (zll_main_multiply1792_inR21[128:1], zll_main_multiply1792_inR21[0], zll_main_multiply1792_outR21);
  assign zll_main_multiply1788_inR12 = {zll_main_multiply1411_in[256:129], zll_main_multiply1411_in[128:1], zll_main_multiply1411_in[0]};
  ZLL_Main_multiply1788  instR85 (zll_main_multiply1788_inR12[256:129], zll_main_multiply1788_inR12[128:1], zll_main_multiply1788_outR12);
  assign zll_main_multiply101_in = {zll_main_multiply138_in[383:256], zll_main_multiply138_in[127:0], (zll_main_multiply1788_inR12[0] == 1'h1) ? zll_main_multiply1788_outR12 : zll_main_multiply1792_outR21};
  assign id_inR65 = zll_main_multiply101_in[255:128];
  assign rewire_prelude_not_inR21 = id_inR65[0];
  ReWire_Prelude_not  instR86 (rewire_prelude_not_inR21[0], rewire_prelude_not_outR21);
  assign zll_main_multiply1785_inR21 = {zll_main_multiply101_in[255:128], rewire_prelude_not_outR21};
  ZLL_Main_multiply1785  instR87 (zll_main_multiply1785_inR21[128:1], zll_main_multiply1785_inR21[0], zll_main_multiply1785_outR21);
  assign zll_main_multiply686_in = {zll_main_multiply101_in[127:0], zll_main_multiply101_in[383:256], zll_main_multiply1785_outR21};
  assign id_inR66 = zll_main_multiply686_in[255:128];
  assign zll_main_multiply1013_in = {zll_main_multiply686_in[127:0], zll_main_multiply686_in[383:256], zll_main_multiply686_in[255:128], id_inR66[105]};
  assign id_inR67 = zll_main_multiply1013_in[128:1];
  assign zll_main_multiply1792_inR22 = {zll_main_multiply1013_in[256:129], id_inR67[105]};
  ZLL_Main_multiply1792  instR88 (zll_main_multiply1792_inR22[128:1], zll_main_multiply1792_inR22[0], zll_main_multiply1792_outR22);
  assign zll_main_multiply1788_inR13 = {zll_main_multiply1013_in[384:257], zll_main_multiply1013_in[256:129], zll_main_multiply1013_in[0]};
  ZLL_Main_multiply1788  instR89 (zll_main_multiply1788_inR13[256:129], zll_main_multiply1788_inR13[128:1], zll_main_multiply1788_outR13);
  assign zll_main_multiply1487_in = {zll_main_multiply686_in[127:0], zll_main_multiply686_in[255:128], (zll_main_multiply1788_inR13[0] == 1'h1) ? zll_main_multiply1788_outR13 : zll_main_multiply1792_outR22};
  assign id_inR68 = zll_main_multiply1487_in[383:256];
  assign rewire_prelude_not_inR22 = id_inR68[0];
  ReWire_Prelude_not  instR90 (rewire_prelude_not_inR22[0], rewire_prelude_not_outR22);
  assign zll_main_multiply1785_inR22 = {zll_main_multiply1487_in[383:256], rewire_prelude_not_outR22};
  ZLL_Main_multiply1785  instR91 (zll_main_multiply1785_inR22[128:1], zll_main_multiply1785_inR22[0], zll_main_multiply1785_outR22);
  assign zll_main_multiply178_in = {zll_main_multiply1487_in[127:0], zll_main_multiply1487_in[255:128], zll_main_multiply1785_outR22};
  assign id_inR69 = zll_main_multiply178_in[255:128];
  assign zll_main_multiply952_in = {zll_main_multiply178_in[383:256], zll_main_multiply178_in[127:0], zll_main_multiply178_in[255:128], id_inR69[104]};
  assign id_inR70 = zll_main_multiply952_in[128:1];
  assign zll_main_multiply1792_inR23 = {zll_main_multiply952_in[384:257], id_inR70[104]};
  ZLL_Main_multiply1792  instR92 (zll_main_multiply1792_inR23[128:1], zll_main_multiply1792_inR23[0], zll_main_multiply1792_outR23);
  assign zll_main_multiply1749_inR9 = {zll_main_multiply952_in[384:257], zll_main_multiply952_in[256:129], zll_main_multiply952_in[0]};
  ZLL_Main_multiply1749  instR93 (zll_main_multiply1749_inR9[256:129], zll_main_multiply1749_inR9[128:1], zll_main_multiply1749_outR9);
  assign zll_main_multiply148_in = {zll_main_multiply178_in[127:0], zll_main_multiply178_in[255:128], (zll_main_multiply1749_inR9[0] == 1'h1) ? zll_main_multiply1749_outR9 : zll_main_multiply1792_outR23};
  assign id_inR71 = zll_main_multiply148_in[383:256];
  assign rewire_prelude_not_inR23 = id_inR71[0];
  ReWire_Prelude_not  instR94 (rewire_prelude_not_inR23[0], rewire_prelude_not_outR23);
  assign zll_main_multiply1785_inR23 = {zll_main_multiply148_in[383:256], rewire_prelude_not_outR23};
  ZLL_Main_multiply1785  instR95 (zll_main_multiply1785_inR23[128:1], zll_main_multiply1785_inR23[0], zll_main_multiply1785_outR23);
  assign zll_main_multiply485_in = {zll_main_multiply148_in[255:128], zll_main_multiply148_in[127:0], zll_main_multiply1785_outR23};
  assign id_inR72 = zll_main_multiply485_in[383:256];
  assign zll_main_multiply1592_in = {zll_main_multiply485_in[127:0], zll_main_multiply485_in[383:256], zll_main_multiply485_in[255:128], id_inR72[103]};
  assign id_inR73 = zll_main_multiply1592_in[256:129];
  assign zll_main_multiply1792_inR24 = {zll_main_multiply1592_in[128:1], id_inR73[103]};
  ZLL_Main_multiply1792  instR96 (zll_main_multiply1792_inR24[128:1], zll_main_multiply1792_inR24[0], zll_main_multiply1792_outR24);
  assign zll_main_multiply1788_inR14 = {zll_main_multiply1592_in[384:257], zll_main_multiply1592_in[128:1], zll_main_multiply1592_in[0]};
  ZLL_Main_multiply1788  instR97 (zll_main_multiply1788_inR14[256:129], zll_main_multiply1788_inR14[128:1], zll_main_multiply1788_outR14);
  assign zll_main_multiply879_in = {zll_main_multiply485_in[127:0], zll_main_multiply485_in[383:256], (zll_main_multiply1788_inR14[0] == 1'h1) ? zll_main_multiply1788_outR14 : zll_main_multiply1792_outR24};
  assign id_inR74 = zll_main_multiply879_in[383:256];
  assign rewire_prelude_not_inR24 = id_inR74[0];
  ReWire_Prelude_not  instR98 (rewire_prelude_not_inR24[0], rewire_prelude_not_outR24);
  assign zll_main_multiply1785_inR24 = {zll_main_multiply879_in[383:256], rewire_prelude_not_outR24};
  ZLL_Main_multiply1785  instR99 (zll_main_multiply1785_inR24[128:1], zll_main_multiply1785_inR24[0], zll_main_multiply1785_outR24);
  assign zll_main_multiply1327_in = {zll_main_multiply879_in[127:0], zll_main_multiply879_in[255:128], zll_main_multiply1785_outR24};
  assign id_inR75 = zll_main_multiply1327_in[255:128];
  assign zll_main_multiply724_in = {zll_main_multiply1327_in[383:256], zll_main_multiply1327_in[255:128], zll_main_multiply1327_in[127:0], id_inR75[102]};
  assign id_inR76 = zll_main_multiply724_in[256:129];
  assign zll_main_multiply1792_inR25 = {zll_main_multiply724_in[384:257], id_inR76[102]};
  ZLL_Main_multiply1792  instR100 (zll_main_multiply1792_inR25[128:1], zll_main_multiply1792_inR25[0], zll_main_multiply1792_outR25);
  assign zll_main_multiply1749_inR10 = {zll_main_multiply724_in[384:257], zll_main_multiply724_in[128:1], zll_main_multiply724_in[0]};
  ZLL_Main_multiply1749  instR101 (zll_main_multiply1749_inR10[256:129], zll_main_multiply1749_inR10[128:1], zll_main_multiply1749_outR10);
  assign zll_main_multiply904_in = {zll_main_multiply1327_in[255:128], zll_main_multiply1327_in[127:0], (zll_main_multiply1749_inR10[0] == 1'h1) ? zll_main_multiply1749_outR10 : zll_main_multiply1792_outR25};
  assign id_inR77 = zll_main_multiply904_in[255:128];
  assign rewire_prelude_not_inR25 = id_inR77[0];
  ReWire_Prelude_not  instR102 (rewire_prelude_not_inR25[0], rewire_prelude_not_outR25);
  assign zll_main_multiply1785_inR25 = {zll_main_multiply904_in[255:128], rewire_prelude_not_outR25};
  ZLL_Main_multiply1785  instR103 (zll_main_multiply1785_inR25[128:1], zll_main_multiply1785_inR25[0], zll_main_multiply1785_outR25);
  assign zll_main_multiply705_in = {zll_main_multiply904_in[127:0], zll_main_multiply904_in[383:256], zll_main_multiply1785_outR25};
  assign id_inR78 = zll_main_multiply705_in[255:128];
  assign zll_main_multiply627_in = {zll_main_multiply705_in[127:0], zll_main_multiply705_in[383:256], zll_main_multiply705_in[255:128], id_inR78[101]};
  assign id_inR79 = zll_main_multiply627_in[128:1];
  assign zll_main_multiply1792_inR26 = {zll_main_multiply627_in[256:129], id_inR79[101]};
  ZLL_Main_multiply1792  instR104 (zll_main_multiply1792_inR26[128:1], zll_main_multiply1792_inR26[0], zll_main_multiply1792_outR26);
  assign zll_main_multiply1788_inR15 = {zll_main_multiply627_in[384:257], zll_main_multiply627_in[256:129], zll_main_multiply627_in[0]};
  ZLL_Main_multiply1788  instR105 (zll_main_multiply1788_inR15[256:129], zll_main_multiply1788_inR15[128:1], zll_main_multiply1788_outR15);
  assign zll_main_multiply847_in = {zll_main_multiply705_in[127:0], zll_main_multiply705_in[255:128], (zll_main_multiply1788_inR15[0] == 1'h1) ? zll_main_multiply1788_outR15 : zll_main_multiply1792_outR26};
  assign id_inR80 = zll_main_multiply847_in[383:256];
  assign rewire_prelude_not_inR26 = id_inR80[0];
  ReWire_Prelude_not  instR106 (rewire_prelude_not_inR26[0], rewire_prelude_not_outR26);
  assign zll_main_multiply1785_inR26 = {zll_main_multiply847_in[383:256], rewire_prelude_not_outR26};
  ZLL_Main_multiply1785  instR107 (zll_main_multiply1785_inR26[128:1], zll_main_multiply1785_inR26[0], zll_main_multiply1785_outR26);
  assign zll_main_multiply560_in = {zll_main_multiply847_in[127:0], zll_main_multiply847_in[255:128], zll_main_multiply1785_outR26};
  assign id_inR81 = zll_main_multiply560_in[255:128];
  assign zll_main_multiply901_in = {zll_main_multiply560_in[127:0], zll_main_multiply560_in[383:256], zll_main_multiply560_in[255:128], id_inR81[100]};
  assign id_inR82 = zll_main_multiply901_in[128:1];
  assign zll_main_multiply1792_inR27 = {zll_main_multiply901_in[256:129], id_inR82[100]};
  ZLL_Main_multiply1792  instR108 (zll_main_multiply1792_inR27[128:1], zll_main_multiply1792_inR27[0], zll_main_multiply1792_outR27);
  assign zll_main_multiply1788_inR16 = {zll_main_multiply901_in[384:257], zll_main_multiply901_in[256:129], zll_main_multiply901_in[0]};
  ZLL_Main_multiply1788  instR109 (zll_main_multiply1788_inR16[256:129], zll_main_multiply1788_inR16[128:1], zll_main_multiply1788_outR16);
  assign zll_main_multiply420_in = {zll_main_multiply560_in[127:0], zll_main_multiply560_in[255:128], (zll_main_multiply1788_inR16[0] == 1'h1) ? zll_main_multiply1788_outR16 : zll_main_multiply1792_outR27};
  assign id_inR83 = zll_main_multiply420_in[383:256];
  assign rewire_prelude_not_inR27 = id_inR83[0];
  ReWire_Prelude_not  instR110 (rewire_prelude_not_inR27[0], rewire_prelude_not_outR27);
  assign zll_main_multiply1785_inR27 = {zll_main_multiply420_in[383:256], rewire_prelude_not_outR27};
  ZLL_Main_multiply1785  instR111 (zll_main_multiply1785_inR27[128:1], zll_main_multiply1785_inR27[0], zll_main_multiply1785_outR27);
  assign zll_main_multiply291_in = {zll_main_multiply420_in[127:0], zll_main_multiply420_in[255:128], zll_main_multiply1785_outR27};
  assign id_inR84 = zll_main_multiply291_in[255:128];
  assign zll_main_multiply185_in = {zll_main_multiply291_in[127:0], zll_main_multiply291_in[383:256], zll_main_multiply291_in[255:128], id_inR84[99]};
  assign id_inR85 = zll_main_multiply185_in[128:1];
  assign zll_main_multiply1792_inR28 = {zll_main_multiply185_in[256:129], id_inR85[99]};
  ZLL_Main_multiply1792  instR112 (zll_main_multiply1792_inR28[128:1], zll_main_multiply1792_inR28[0], zll_main_multiply1792_outR28);
  assign zll_main_multiply1788_inR17 = {zll_main_multiply185_in[384:257], zll_main_multiply185_in[256:129], zll_main_multiply185_in[0]};
  ZLL_Main_multiply1788  instR113 (zll_main_multiply1788_inR17[256:129], zll_main_multiply1788_inR17[128:1], zll_main_multiply1788_outR17);
  assign zll_main_multiply749_in = {zll_main_multiply291_in[127:0], zll_main_multiply291_in[255:128], (zll_main_multiply1788_inR17[0] == 1'h1) ? zll_main_multiply1788_outR17 : zll_main_multiply1792_outR28};
  assign id_inR86 = zll_main_multiply749_in[383:256];
  assign rewire_prelude_not_inR28 = id_inR86[0];
  ReWire_Prelude_not  instR114 (rewire_prelude_not_inR28[0], rewire_prelude_not_outR28);
  assign zll_main_multiply1785_inR28 = {zll_main_multiply749_in[383:256], rewire_prelude_not_outR28};
  ZLL_Main_multiply1785  instR115 (zll_main_multiply1785_inR28[128:1], zll_main_multiply1785_inR28[0], zll_main_multiply1785_outR28);
  assign zll_main_multiply810_in = {zll_main_multiply749_in[255:128], zll_main_multiply749_in[127:0], zll_main_multiply1785_outR28};
  assign id_inR87 = zll_main_multiply810_in[383:256];
  assign zll_main_multiply154_in = {zll_main_multiply810_in[383:256], zll_main_multiply810_in[255:128], zll_main_multiply810_in[127:0], id_inR87[98]};
  assign id_inR88 = zll_main_multiply154_in[384:257];
  assign zll_main_multiply1792_inR29 = {zll_main_multiply154_in[256:129], id_inR88[98]};
  ZLL_Main_multiply1792  instR116 (zll_main_multiply1792_inR29[128:1], zll_main_multiply1792_inR29[0], zll_main_multiply1792_outR29);
  assign zll_main_multiply1749_inR11 = {zll_main_multiply154_in[256:129], zll_main_multiply154_in[128:1], zll_main_multiply154_in[0]};
  ZLL_Main_multiply1749  instR117 (zll_main_multiply1749_inR11[256:129], zll_main_multiply1749_inR11[128:1], zll_main_multiply1749_outR11);
  assign zll_main_multiply1542_in = {zll_main_multiply810_in[383:256], zll_main_multiply810_in[127:0], (zll_main_multiply1749_inR11[0] == 1'h1) ? zll_main_multiply1749_outR11 : zll_main_multiply1792_outR29};
  assign id_inR89 = zll_main_multiply1542_in[255:128];
  assign rewire_prelude_not_inR29 = id_inR89[0];
  ReWire_Prelude_not  instR118 (rewire_prelude_not_inR29[0], rewire_prelude_not_outR29);
  assign zll_main_multiply1785_inR29 = {zll_main_multiply1542_in[255:128], rewire_prelude_not_outR29};
  ZLL_Main_multiply1785  instR119 (zll_main_multiply1785_inR29[128:1], zll_main_multiply1785_inR29[0], zll_main_multiply1785_outR29);
  assign zll_main_multiply1173_in = {zll_main_multiply1542_in[383:256], zll_main_multiply1542_in[127:0], zll_main_multiply1785_outR29};
  assign id_inR90 = zll_main_multiply1173_in[383:256];
  assign zll_main_multiply512_in = {zll_main_multiply1173_in[127:0], zll_main_multiply1173_in[383:256], zll_main_multiply1173_in[255:128], id_inR90[97]};
  assign id_inR91 = zll_main_multiply512_in[256:129];
  assign zll_main_multiply1792_inR30 = {zll_main_multiply512_in[128:1], id_inR91[97]};
  ZLL_Main_multiply1792  instR120 (zll_main_multiply1792_inR30[128:1], zll_main_multiply1792_inR30[0], zll_main_multiply1792_outR30);
  assign zll_main_multiply1788_inR18 = {zll_main_multiply512_in[384:257], zll_main_multiply512_in[128:1], zll_main_multiply512_in[0]};
  ZLL_Main_multiply1788  instR121 (zll_main_multiply1788_inR18[256:129], zll_main_multiply1788_inR18[128:1], zll_main_multiply1788_outR18);
  assign zll_main_multiply66_in = {zll_main_multiply1173_in[127:0], zll_main_multiply1173_in[383:256], (zll_main_multiply1788_inR18[0] == 1'h1) ? zll_main_multiply1788_outR18 : zll_main_multiply1792_outR30};
  assign id_inR92 = zll_main_multiply66_in[383:256];
  assign rewire_prelude_not_inR30 = id_inR92[0];
  ReWire_Prelude_not  instR122 (rewire_prelude_not_inR30[0], rewire_prelude_not_outR30);
  assign zll_main_multiply1785_inR30 = {zll_main_multiply66_in[383:256], rewire_prelude_not_outR30};
  ZLL_Main_multiply1785  instR123 (zll_main_multiply1785_inR30[128:1], zll_main_multiply1785_inR30[0], zll_main_multiply1785_outR30);
  assign zll_main_multiply1574_in = {zll_main_multiply66_in[255:128], zll_main_multiply66_in[127:0], zll_main_multiply1785_outR30};
  assign id_inR93 = zll_main_multiply1574_in[383:256];
  assign zll_main_multiply550_in = {zll_main_multiply1574_in[127:0], zll_main_multiply1574_in[383:256], zll_main_multiply1574_in[255:128], id_inR93[96]};
  assign id_inR94 = zll_main_multiply550_in[256:129];
  assign zll_main_multiply1792_inR31 = {zll_main_multiply550_in[128:1], id_inR94[96]};
  ZLL_Main_multiply1792  instR124 (zll_main_multiply1792_inR31[128:1], zll_main_multiply1792_inR31[0], zll_main_multiply1792_outR31);
  assign zll_main_multiply1788_inR19 = {zll_main_multiply550_in[384:257], zll_main_multiply550_in[128:1], zll_main_multiply550_in[0]};
  ZLL_Main_multiply1788  instR125 (zll_main_multiply1788_inR19[256:129], zll_main_multiply1788_inR19[128:1], zll_main_multiply1788_outR19);
  assign zll_main_multiply1392_in = {zll_main_multiply1574_in[127:0], zll_main_multiply1574_in[383:256], (zll_main_multiply1788_inR19[0] == 1'h1) ? zll_main_multiply1788_outR19 : zll_main_multiply1792_outR31};
  assign id_inR95 = zll_main_multiply1392_in[383:256];
  assign rewire_prelude_not_inR31 = id_inR95[0];
  ReWire_Prelude_not  instR126 (rewire_prelude_not_inR31[0], rewire_prelude_not_outR31);
  assign zll_main_multiply1785_inR31 = {zll_main_multiply1392_in[383:256], rewire_prelude_not_outR31};
  ZLL_Main_multiply1785  instR127 (zll_main_multiply1785_inR31[128:1], zll_main_multiply1785_inR31[0], zll_main_multiply1785_outR31);
  assign zll_main_multiply450_in = {zll_main_multiply1392_in[127:0], zll_main_multiply1392_in[255:128], zll_main_multiply1785_outR31};
  assign id_inR96 = zll_main_multiply450_in[255:128];
  assign zll_main_multiply193_in = {zll_main_multiply450_in[127:0], zll_main_multiply450_in[383:256], zll_main_multiply450_in[255:128], id_inR96[95]};
  assign id_inR97 = zll_main_multiply193_in[128:1];
  assign zll_main_multiply1792_inR32 = {zll_main_multiply193_in[256:129], id_inR97[95]};
  ZLL_Main_multiply1792  instR128 (zll_main_multiply1792_inR32[128:1], zll_main_multiply1792_inR32[0], zll_main_multiply1792_outR32);
  assign zll_main_multiply1788_inR20 = {zll_main_multiply193_in[384:257], zll_main_multiply193_in[256:129], zll_main_multiply193_in[0]};
  ZLL_Main_multiply1788  instR129 (zll_main_multiply1788_inR20[256:129], zll_main_multiply1788_inR20[128:1], zll_main_multiply1788_outR20);
  assign zll_main_multiply633_in = {zll_main_multiply450_in[127:0], zll_main_multiply450_in[255:128], (zll_main_multiply1788_inR20[0] == 1'h1) ? zll_main_multiply1788_outR20 : zll_main_multiply1792_outR32};
  assign id_inR98 = zll_main_multiply633_in[383:256];
  assign rewire_prelude_not_inR32 = id_inR98[0];
  ReWire_Prelude_not  instR130 (rewire_prelude_not_inR32[0], rewire_prelude_not_outR32);
  assign zll_main_multiply1785_inR32 = {zll_main_multiply633_in[383:256], rewire_prelude_not_outR32};
  ZLL_Main_multiply1785  instR131 (zll_main_multiply1785_inR32[128:1], zll_main_multiply1785_inR32[0], zll_main_multiply1785_outR32);
  assign zll_main_multiply1596_in = {zll_main_multiply633_in[127:0], zll_main_multiply633_in[255:128], zll_main_multiply1785_outR32};
  assign id_inR99 = zll_main_multiply1596_in[255:128];
  assign zll_main_multiply315_in = {zll_main_multiply1596_in[383:256], zll_main_multiply1596_in[127:0], zll_main_multiply1596_in[255:128], id_inR99[94]};
  assign id_inR100 = zll_main_multiply315_in[128:1];
  assign zll_main_multiply1792_inR33 = {zll_main_multiply315_in[384:257], id_inR100[94]};
  ZLL_Main_multiply1792  instR132 (zll_main_multiply1792_inR33[128:1], zll_main_multiply1792_inR33[0], zll_main_multiply1792_outR33);
  assign zll_main_multiply1749_inR12 = {zll_main_multiply315_in[384:257], zll_main_multiply315_in[256:129], zll_main_multiply315_in[0]};
  ZLL_Main_multiply1749  instR133 (zll_main_multiply1749_inR12[256:129], zll_main_multiply1749_inR12[128:1], zll_main_multiply1749_outR12);
  assign zll_main_multiply165_in = {zll_main_multiply1596_in[127:0], zll_main_multiply1596_in[255:128], (zll_main_multiply1749_inR12[0] == 1'h1) ? zll_main_multiply1749_outR12 : zll_main_multiply1792_outR33};
  assign id_inR101 = zll_main_multiply165_in[383:256];
  assign rewire_prelude_not_inR33 = id_inR101[0];
  ReWire_Prelude_not  instR134 (rewire_prelude_not_inR33[0], rewire_prelude_not_outR33);
  assign zll_main_multiply1785_inR33 = {zll_main_multiply165_in[383:256], rewire_prelude_not_outR33};
  ZLL_Main_multiply1785  instR135 (zll_main_multiply1785_inR33[128:1], zll_main_multiply1785_inR33[0], zll_main_multiply1785_outR33);
  assign zll_main_multiply934_in = {zll_main_multiply165_in[255:128], zll_main_multiply165_in[127:0], zll_main_multiply1785_outR33};
  assign id_inR102 = zll_main_multiply934_in[383:256];
  assign zll_main_multiply738_in = {zll_main_multiply934_in[127:0], zll_main_multiply934_in[383:256], zll_main_multiply934_in[255:128], id_inR102[93]};
  assign id_inR103 = zll_main_multiply738_in[256:129];
  assign zll_main_multiply1792_inR34 = {zll_main_multiply738_in[128:1], id_inR103[93]};
  ZLL_Main_multiply1792  instR136 (zll_main_multiply1792_inR34[128:1], zll_main_multiply1792_inR34[0], zll_main_multiply1792_outR34);
  assign zll_main_multiply1788_inR21 = {zll_main_multiply738_in[384:257], zll_main_multiply738_in[128:1], zll_main_multiply738_in[0]};
  ZLL_Main_multiply1788  instR137 (zll_main_multiply1788_inR21[256:129], zll_main_multiply1788_inR21[128:1], zll_main_multiply1788_outR21);
  assign zll_main_multiply278_in = {zll_main_multiply934_in[127:0], zll_main_multiply934_in[383:256], (zll_main_multiply1788_inR21[0] == 1'h1) ? zll_main_multiply1788_outR21 : zll_main_multiply1792_outR34};
  assign id_inR104 = zll_main_multiply278_in[383:256];
  assign rewire_prelude_not_inR34 = id_inR104[0];
  ReWire_Prelude_not  instR138 (rewire_prelude_not_inR34[0], rewire_prelude_not_outR34);
  assign zll_main_multiply1785_inR34 = {zll_main_multiply278_in[383:256], rewire_prelude_not_outR34};
  ZLL_Main_multiply1785  instR139 (zll_main_multiply1785_inR34[128:1], zll_main_multiply1785_inR34[0], zll_main_multiply1785_outR34);
  assign zll_main_multiply271_in = {zll_main_multiply278_in[127:0], zll_main_multiply278_in[255:128], zll_main_multiply1785_outR34};
  assign id_inR105 = zll_main_multiply271_in[255:128];
  assign zll_main_multiply1331_in = {zll_main_multiply271_in[127:0], zll_main_multiply271_in[383:256], zll_main_multiply271_in[255:128], id_inR105[92]};
  assign id_inR106 = zll_main_multiply1331_in[128:1];
  assign zll_main_multiply1792_inR35 = {zll_main_multiply1331_in[256:129], id_inR106[92]};
  ZLL_Main_multiply1792  instR140 (zll_main_multiply1792_inR35[128:1], zll_main_multiply1792_inR35[0], zll_main_multiply1792_outR35);
  assign zll_main_multiply1788_inR22 = {zll_main_multiply1331_in[384:257], zll_main_multiply1331_in[256:129], zll_main_multiply1331_in[0]};
  ZLL_Main_multiply1788  instR141 (zll_main_multiply1788_inR22[256:129], zll_main_multiply1788_inR22[128:1], zll_main_multiply1788_outR22);
  assign zll_main_multiply993_in = {zll_main_multiply271_in[127:0], zll_main_multiply271_in[255:128], (zll_main_multiply1788_inR22[0] == 1'h1) ? zll_main_multiply1788_outR22 : zll_main_multiply1792_outR35};
  assign id_inR107 = zll_main_multiply993_in[383:256];
  assign rewire_prelude_not_inR35 = id_inR107[0];
  ReWire_Prelude_not  instR142 (rewire_prelude_not_inR35[0], rewire_prelude_not_outR35);
  assign zll_main_multiply1785_inR35 = {zll_main_multiply993_in[383:256], rewire_prelude_not_outR35};
  ZLL_Main_multiply1785  instR143 (zll_main_multiply1785_inR35[128:1], zll_main_multiply1785_inR35[0], zll_main_multiply1785_outR35);
  assign zll_main_multiply1389_in = {zll_main_multiply993_in[127:0], zll_main_multiply993_in[255:128], zll_main_multiply1785_outR35};
  assign id_inR108 = zll_main_multiply1389_in[255:128];
  assign zll_main_multiply1343_in = {zll_main_multiply1389_in[383:256], zll_main_multiply1389_in[127:0], zll_main_multiply1389_in[255:128], id_inR108[91]};
  assign id_inR109 = zll_main_multiply1343_in[128:1];
  assign zll_main_multiply1792_inR36 = {zll_main_multiply1343_in[384:257], id_inR109[91]};
  ZLL_Main_multiply1792  instR144 (zll_main_multiply1792_inR36[128:1], zll_main_multiply1792_inR36[0], zll_main_multiply1792_outR36);
  assign zll_main_multiply1749_inR13 = {zll_main_multiply1343_in[384:257], zll_main_multiply1343_in[256:129], zll_main_multiply1343_in[0]};
  ZLL_Main_multiply1749  instR145 (zll_main_multiply1749_inR13[256:129], zll_main_multiply1749_inR13[128:1], zll_main_multiply1749_outR13);
  assign zll_main_multiply873_in = {zll_main_multiply1389_in[127:0], zll_main_multiply1389_in[255:128], (zll_main_multiply1749_inR13[0] == 1'h1) ? zll_main_multiply1749_outR13 : zll_main_multiply1792_outR36};
  assign id_inR110 = zll_main_multiply873_in[383:256];
  assign rewire_prelude_not_inR36 = id_inR110[0];
  ReWire_Prelude_not  instR146 (rewire_prelude_not_inR36[0], rewire_prelude_not_outR36);
  assign zll_main_multiply1785_inR36 = {zll_main_multiply873_in[383:256], rewire_prelude_not_outR36};
  ZLL_Main_multiply1785  instR147 (zll_main_multiply1785_inR36[128:1], zll_main_multiply1785_inR36[0], zll_main_multiply1785_outR36);
  assign zll_main_multiply1626_in = {zll_main_multiply873_in[127:0], zll_main_multiply873_in[255:128], zll_main_multiply1785_outR36};
  assign id_inR111 = zll_main_multiply1626_in[255:128];
  assign zll_main_multiply350_in = {zll_main_multiply1626_in[383:256], zll_main_multiply1626_in[127:0], zll_main_multiply1626_in[255:128], id_inR111[90]};
  assign id_inR112 = zll_main_multiply350_in[128:1];
  assign zll_main_multiply1792_inR37 = {zll_main_multiply350_in[384:257], id_inR112[90]};
  ZLL_Main_multiply1792  instR148 (zll_main_multiply1792_inR37[128:1], zll_main_multiply1792_inR37[0], zll_main_multiply1792_outR37);
  assign zll_main_multiply1749_inR14 = {zll_main_multiply350_in[384:257], zll_main_multiply350_in[256:129], zll_main_multiply350_in[0]};
  ZLL_Main_multiply1749  instR149 (zll_main_multiply1749_inR14[256:129], zll_main_multiply1749_inR14[128:1], zll_main_multiply1749_outR14);
  assign zll_main_multiply421_in = {zll_main_multiply1626_in[127:0], zll_main_multiply1626_in[255:128], (zll_main_multiply1749_inR14[0] == 1'h1) ? zll_main_multiply1749_outR14 : zll_main_multiply1792_outR37};
  assign id_inR113 = zll_main_multiply421_in[383:256];
  assign rewire_prelude_not_inR37 = id_inR113[0];
  ReWire_Prelude_not  instR150 (rewire_prelude_not_inR37[0], rewire_prelude_not_outR37);
  assign zll_main_multiply1785_inR37 = {zll_main_multiply421_in[383:256], rewire_prelude_not_outR37};
  ZLL_Main_multiply1785  instR151 (zll_main_multiply1785_inR37[128:1], zll_main_multiply1785_inR37[0], zll_main_multiply1785_outR37);
  assign zll_main_multiply556_in = {zll_main_multiply421_in[127:0], zll_main_multiply421_in[255:128], zll_main_multiply1785_outR37};
  assign id_inR114 = zll_main_multiply556_in[255:128];
  assign zll_main_multiply1036_in = {zll_main_multiply556_in[383:256], zll_main_multiply556_in[255:128], zll_main_multiply556_in[127:0], id_inR114[89]};
  assign id_inR115 = zll_main_multiply1036_in[256:129];
  assign zll_main_multiply1792_inR38 = {zll_main_multiply1036_in[384:257], id_inR115[89]};
  ZLL_Main_multiply1792  instR152 (zll_main_multiply1792_inR38[128:1], zll_main_multiply1792_inR38[0], zll_main_multiply1792_outR38);
  assign zll_main_multiply1749_inR15 = {zll_main_multiply1036_in[384:257], zll_main_multiply1036_in[128:1], zll_main_multiply1036_in[0]};
  ZLL_Main_multiply1749  instR153 (zll_main_multiply1749_inR15[256:129], zll_main_multiply1749_inR15[128:1], zll_main_multiply1749_outR15);
  assign zll_main_multiply22_in = {zll_main_multiply556_in[255:128], zll_main_multiply556_in[127:0], (zll_main_multiply1749_inR15[0] == 1'h1) ? zll_main_multiply1749_outR15 : zll_main_multiply1792_outR38};
  assign id_inR116 = zll_main_multiply22_in[255:128];
  assign rewire_prelude_not_inR38 = id_inR116[0];
  ReWire_Prelude_not  instR154 (rewire_prelude_not_inR38[0], rewire_prelude_not_outR38);
  assign zll_main_multiply1785_inR38 = {zll_main_multiply22_in[255:128], rewire_prelude_not_outR38};
  ZLL_Main_multiply1785  instR155 (zll_main_multiply1785_inR38[128:1], zll_main_multiply1785_inR38[0], zll_main_multiply1785_outR38);
  assign zll_main_multiply905_in = {zll_main_multiply22_in[127:0], zll_main_multiply22_in[383:256], zll_main_multiply1785_outR38};
  assign id_inR117 = zll_main_multiply905_in[255:128];
  assign zll_main_multiply1518_in = {zll_main_multiply905_in[383:256], zll_main_multiply905_in[127:0], zll_main_multiply905_in[255:128], id_inR117[88]};
  assign id_inR118 = zll_main_multiply1518_in[128:1];
  assign zll_main_multiply1792_inR39 = {zll_main_multiply1518_in[384:257], id_inR118[88]};
  ZLL_Main_multiply1792  instR156 (zll_main_multiply1792_inR39[128:1], zll_main_multiply1792_inR39[0], zll_main_multiply1792_outR39);
  assign zll_main_multiply1749_inR16 = {zll_main_multiply1518_in[384:257], zll_main_multiply1518_in[256:129], zll_main_multiply1518_in[0]};
  ZLL_Main_multiply1749  instR157 (zll_main_multiply1749_inR16[256:129], zll_main_multiply1749_inR16[128:1], zll_main_multiply1749_outR16);
  assign zll_main_multiply403_in = {zll_main_multiply905_in[127:0], zll_main_multiply905_in[255:128], (zll_main_multiply1749_inR16[0] == 1'h1) ? zll_main_multiply1749_outR16 : zll_main_multiply1792_outR39};
  assign id_inR119 = zll_main_multiply403_in[383:256];
  assign rewire_prelude_not_inR39 = id_inR119[0];
  ReWire_Prelude_not  instR158 (rewire_prelude_not_inR39[0], rewire_prelude_not_outR39);
  assign zll_main_multiply1785_inR39 = {zll_main_multiply403_in[383:256], rewire_prelude_not_outR39};
  ZLL_Main_multiply1785  instR159 (zll_main_multiply1785_inR39[128:1], zll_main_multiply1785_inR39[0], zll_main_multiply1785_outR39);
  assign zll_main_multiply644_in = {zll_main_multiply403_in[127:0], zll_main_multiply403_in[255:128], zll_main_multiply1785_outR39};
  assign id_inR120 = zll_main_multiply644_in[255:128];
  assign zll_main_multiply431_in = {zll_main_multiply644_in[383:256], zll_main_multiply644_in[255:128], zll_main_multiply644_in[127:0], id_inR120[87]};
  assign id_inR121 = zll_main_multiply431_in[256:129];
  assign zll_main_multiply1792_inR40 = {zll_main_multiply431_in[384:257], id_inR121[87]};
  ZLL_Main_multiply1792  instR160 (zll_main_multiply1792_inR40[128:1], zll_main_multiply1792_inR40[0], zll_main_multiply1792_outR40);
  assign zll_main_multiply1749_inR17 = {zll_main_multiply431_in[384:257], zll_main_multiply431_in[128:1], zll_main_multiply431_in[0]};
  ZLL_Main_multiply1749  instR161 (zll_main_multiply1749_inR17[256:129], zll_main_multiply1749_inR17[128:1], zll_main_multiply1749_outR17);
  assign zll_main_multiply256_in = {zll_main_multiply644_in[255:128], zll_main_multiply644_in[127:0], (zll_main_multiply1749_inR17[0] == 1'h1) ? zll_main_multiply1749_outR17 : zll_main_multiply1792_outR40};
  assign id_inR122 = zll_main_multiply256_in[255:128];
  assign rewire_prelude_not_inR40 = id_inR122[0];
  ReWire_Prelude_not  instR162 (rewire_prelude_not_inR40[0], rewire_prelude_not_outR40);
  assign zll_main_multiply1785_inR40 = {zll_main_multiply256_in[255:128], rewire_prelude_not_outR40};
  ZLL_Main_multiply1785  instR163 (zll_main_multiply1785_inR40[128:1], zll_main_multiply1785_inR40[0], zll_main_multiply1785_outR40);
  assign zll_main_multiply198_in = {zll_main_multiply256_in[383:256], zll_main_multiply256_in[127:0], zll_main_multiply1785_outR40};
  assign id_inR123 = zll_main_multiply198_in[383:256];
  assign zll_main_multiply846_in = {zll_main_multiply198_in[383:256], zll_main_multiply198_in[255:128], zll_main_multiply198_in[127:0], id_inR123[86]};
  assign id_inR124 = zll_main_multiply846_in[384:257];
  assign zll_main_multiply1792_inR41 = {zll_main_multiply846_in[256:129], id_inR124[86]};
  ZLL_Main_multiply1792  instR164 (zll_main_multiply1792_inR41[128:1], zll_main_multiply1792_inR41[0], zll_main_multiply1792_outR41);
  assign zll_main_multiply1749_inR18 = {zll_main_multiply846_in[256:129], zll_main_multiply846_in[128:1], zll_main_multiply846_in[0]};
  ZLL_Main_multiply1749  instR165 (zll_main_multiply1749_inR18[256:129], zll_main_multiply1749_inR18[128:1], zll_main_multiply1749_outR18);
  assign zll_main_multiply25_in = {zll_main_multiply198_in[383:256], zll_main_multiply198_in[127:0], (zll_main_multiply1749_inR18[0] == 1'h1) ? zll_main_multiply1749_outR18 : zll_main_multiply1792_outR41};
  assign id_inR125 = zll_main_multiply25_in[255:128];
  assign rewire_prelude_not_inR41 = id_inR125[0];
  ReWire_Prelude_not  instR166 (rewire_prelude_not_inR41[0], rewire_prelude_not_outR41);
  assign zll_main_multiply1785_inR41 = {zll_main_multiply25_in[255:128], rewire_prelude_not_outR41};
  ZLL_Main_multiply1785  instR167 (zll_main_multiply1785_inR41[128:1], zll_main_multiply1785_inR41[0], zll_main_multiply1785_outR41);
  assign zll_main_multiply381_in = {zll_main_multiply25_in[383:256], zll_main_multiply25_in[127:0], zll_main_multiply1785_outR41};
  assign id_inR126 = zll_main_multiply381_in[383:256];
  assign zll_main_multiply285_in = {zll_main_multiply381_in[127:0], zll_main_multiply381_in[383:256], zll_main_multiply381_in[255:128], id_inR126[85]};
  assign id_inR127 = zll_main_multiply285_in[256:129];
  assign zll_main_multiply1792_inR42 = {zll_main_multiply285_in[128:1], id_inR127[85]};
  ZLL_Main_multiply1792  instR168 (zll_main_multiply1792_inR42[128:1], zll_main_multiply1792_inR42[0], zll_main_multiply1792_outR42);
  assign zll_main_multiply1788_inR23 = {zll_main_multiply285_in[384:257], zll_main_multiply285_in[128:1], zll_main_multiply285_in[0]};
  ZLL_Main_multiply1788  instR169 (zll_main_multiply1788_inR23[256:129], zll_main_multiply1788_inR23[128:1], zll_main_multiply1788_outR23);
  assign zll_main_multiply1355_in = {zll_main_multiply381_in[127:0], zll_main_multiply381_in[383:256], (zll_main_multiply1788_inR23[0] == 1'h1) ? zll_main_multiply1788_outR23 : zll_main_multiply1792_outR42};
  assign id_inR128 = zll_main_multiply1355_in[383:256];
  assign rewire_prelude_not_inR42 = id_inR128[0];
  ReWire_Prelude_not  instR170 (rewire_prelude_not_inR42[0], rewire_prelude_not_outR42);
  assign zll_main_multiply1785_inR42 = {zll_main_multiply1355_in[383:256], rewire_prelude_not_outR42};
  ZLL_Main_multiply1785  instR171 (zll_main_multiply1785_inR42[128:1], zll_main_multiply1785_inR42[0], zll_main_multiply1785_outR42);
  assign zll_main_multiply1141_in = {zll_main_multiply1355_in[127:0], zll_main_multiply1355_in[255:128], zll_main_multiply1785_outR42};
  assign id_inR129 = zll_main_multiply1141_in[255:128];
  assign zll_main_multiply188_in = {zll_main_multiply1141_in[127:0], zll_main_multiply1141_in[383:256], zll_main_multiply1141_in[255:128], id_inR129[84]};
  assign id_inR130 = zll_main_multiply188_in[128:1];
  assign zll_main_multiply1792_inR43 = {zll_main_multiply188_in[256:129], id_inR130[84]};
  ZLL_Main_multiply1792  instR172 (zll_main_multiply1792_inR43[128:1], zll_main_multiply1792_inR43[0], zll_main_multiply1792_outR43);
  assign zll_main_multiply1788_inR24 = {zll_main_multiply188_in[384:257], zll_main_multiply188_in[256:129], zll_main_multiply188_in[0]};
  ZLL_Main_multiply1788  instR173 (zll_main_multiply1788_inR24[256:129], zll_main_multiply1788_inR24[128:1], zll_main_multiply1788_outR24);
  assign zll_main_multiply558_in = {zll_main_multiply1141_in[127:0], zll_main_multiply1141_in[255:128], (zll_main_multiply1788_inR24[0] == 1'h1) ? zll_main_multiply1788_outR24 : zll_main_multiply1792_outR43};
  assign id_inR131 = zll_main_multiply558_in[383:256];
  assign rewire_prelude_not_inR43 = id_inR131[0];
  ReWire_Prelude_not  instR174 (rewire_prelude_not_inR43[0], rewire_prelude_not_outR43);
  assign zll_main_multiply1785_inR43 = {zll_main_multiply558_in[383:256], rewire_prelude_not_outR43};
  ZLL_Main_multiply1785  instR175 (zll_main_multiply1785_inR43[128:1], zll_main_multiply1785_inR43[0], zll_main_multiply1785_outR43);
  assign zll_main_multiply706_in = {zll_main_multiply558_in[255:128], zll_main_multiply558_in[127:0], zll_main_multiply1785_outR43};
  assign id_inR132 = zll_main_multiply706_in[383:256];
  assign zll_main_multiply323_in = {zll_main_multiply706_in[383:256], zll_main_multiply706_in[255:128], zll_main_multiply706_in[127:0], id_inR132[83]};
  assign id_inR133 = zll_main_multiply323_in[384:257];
  assign zll_main_multiply1792_inR44 = {zll_main_multiply323_in[256:129], id_inR133[83]};
  ZLL_Main_multiply1792  instR176 (zll_main_multiply1792_inR44[128:1], zll_main_multiply1792_inR44[0], zll_main_multiply1792_outR44);
  assign zll_main_multiply1749_inR19 = {zll_main_multiply323_in[256:129], zll_main_multiply323_in[128:1], zll_main_multiply323_in[0]};
  ZLL_Main_multiply1749  instR177 (zll_main_multiply1749_inR19[256:129], zll_main_multiply1749_inR19[128:1], zll_main_multiply1749_outR19);
  assign zll_main_multiply1675_in = {zll_main_multiply706_in[383:256], zll_main_multiply706_in[127:0], (zll_main_multiply1749_inR19[0] == 1'h1) ? zll_main_multiply1749_outR19 : zll_main_multiply1792_outR44};
  assign id_inR134 = zll_main_multiply1675_in[255:128];
  assign rewire_prelude_not_inR44 = id_inR134[0];
  ReWire_Prelude_not  instR178 (rewire_prelude_not_inR44[0], rewire_prelude_not_outR44);
  assign zll_main_multiply1785_inR44 = {zll_main_multiply1675_in[255:128], rewire_prelude_not_outR44};
  ZLL_Main_multiply1785  instR179 (zll_main_multiply1785_inR44[128:1], zll_main_multiply1785_inR44[0], zll_main_multiply1785_outR44);
  assign zll_main_multiply863_in = {zll_main_multiply1675_in[127:0], zll_main_multiply1675_in[383:256], zll_main_multiply1785_outR44};
  assign id_inR135 = zll_main_multiply863_in[255:128];
  assign zll_main_multiply1246_in = {zll_main_multiply863_in[383:256], zll_main_multiply863_in[255:128], zll_main_multiply863_in[127:0], id_inR135[82]};
  assign id_inR136 = zll_main_multiply1246_in[256:129];
  assign zll_main_multiply1792_inR45 = {zll_main_multiply1246_in[384:257], id_inR136[82]};
  ZLL_Main_multiply1792  instR180 (zll_main_multiply1792_inR45[128:1], zll_main_multiply1792_inR45[0], zll_main_multiply1792_outR45);
  assign zll_main_multiply1749_inR20 = {zll_main_multiply1246_in[384:257], zll_main_multiply1246_in[128:1], zll_main_multiply1246_in[0]};
  ZLL_Main_multiply1749  instR181 (zll_main_multiply1749_inR20[256:129], zll_main_multiply1749_inR20[128:1], zll_main_multiply1749_outR20);
  assign zll_main_multiply190_in = {zll_main_multiply863_in[255:128], zll_main_multiply863_in[127:0], (zll_main_multiply1749_inR20[0] == 1'h1) ? zll_main_multiply1749_outR20 : zll_main_multiply1792_outR45};
  assign id_inR137 = zll_main_multiply190_in[255:128];
  assign rewire_prelude_not_inR45 = id_inR137[0];
  ReWire_Prelude_not  instR182 (rewire_prelude_not_inR45[0], rewire_prelude_not_outR45);
  assign zll_main_multiply1785_inR45 = {zll_main_multiply190_in[255:128], rewire_prelude_not_outR45};
  ZLL_Main_multiply1785  instR183 (zll_main_multiply1785_inR45[128:1], zll_main_multiply1785_inR45[0], zll_main_multiply1785_outR45);
  assign zll_main_multiply7_in = {zll_main_multiply190_in[127:0], zll_main_multiply190_in[383:256], zll_main_multiply1785_outR45};
  assign id_inR138 = zll_main_multiply7_in[255:128];
  assign zll_main_multiply1112_in = {zll_main_multiply7_in[383:256], zll_main_multiply7_in[255:128], zll_main_multiply7_in[127:0], id_inR138[81]};
  assign id_inR139 = zll_main_multiply1112_in[256:129];
  assign zll_main_multiply1792_inR46 = {zll_main_multiply1112_in[384:257], id_inR139[81]};
  ZLL_Main_multiply1792  instR184 (zll_main_multiply1792_inR46[128:1], zll_main_multiply1792_inR46[0], zll_main_multiply1792_outR46);
  assign zll_main_multiply1749_inR21 = {zll_main_multiply1112_in[384:257], zll_main_multiply1112_in[128:1], zll_main_multiply1112_in[0]};
  ZLL_Main_multiply1749  instR185 (zll_main_multiply1749_inR21[256:129], zll_main_multiply1749_inR21[128:1], zll_main_multiply1749_outR21);
  assign zll_main_multiply906_in = {zll_main_multiply7_in[255:128], zll_main_multiply7_in[127:0], (zll_main_multiply1749_inR21[0] == 1'h1) ? zll_main_multiply1749_outR21 : zll_main_multiply1792_outR46};
  assign id_inR140 = zll_main_multiply906_in[255:128];
  assign rewire_prelude_not_inR46 = id_inR140[0];
  ReWire_Prelude_not  instR186 (rewire_prelude_not_inR46[0], rewire_prelude_not_outR46);
  assign zll_main_multiply1785_inR46 = {zll_main_multiply906_in[255:128], rewire_prelude_not_outR46};
  ZLL_Main_multiply1785  instR187 (zll_main_multiply1785_inR46[128:1], zll_main_multiply1785_inR46[0], zll_main_multiply1785_outR46);
  assign zll_main_multiply865_in = {zll_main_multiply906_in[383:256], zll_main_multiply906_in[127:0], zll_main_multiply1785_outR46};
  assign id_inR141 = zll_main_multiply865_in[383:256];
  assign zll_main_multiply1034_in = {zll_main_multiply865_in[127:0], zll_main_multiply865_in[383:256], zll_main_multiply865_in[255:128], id_inR141[80]};
  assign id_inR142 = zll_main_multiply1034_in[256:129];
  assign zll_main_multiply1792_inR47 = {zll_main_multiply1034_in[128:1], id_inR142[80]};
  ZLL_Main_multiply1792  instR188 (zll_main_multiply1792_inR47[128:1], zll_main_multiply1792_inR47[0], zll_main_multiply1792_outR47);
  assign zll_main_multiply1788_inR25 = {zll_main_multiply1034_in[384:257], zll_main_multiply1034_in[128:1], zll_main_multiply1034_in[0]};
  ZLL_Main_multiply1788  instR189 (zll_main_multiply1788_inR25[256:129], zll_main_multiply1788_inR25[128:1], zll_main_multiply1788_outR25);
  assign zll_main_multiply1238_in = {zll_main_multiply865_in[127:0], zll_main_multiply865_in[383:256], (zll_main_multiply1788_inR25[0] == 1'h1) ? zll_main_multiply1788_outR25 : zll_main_multiply1792_outR47};
  assign id_inR143 = zll_main_multiply1238_in[383:256];
  assign rewire_prelude_not_inR47 = id_inR143[0];
  ReWire_Prelude_not  instR190 (rewire_prelude_not_inR47[0], rewire_prelude_not_outR47);
  assign zll_main_multiply1785_inR47 = {zll_main_multiply1238_in[383:256], rewire_prelude_not_outR47};
  ZLL_Main_multiply1785  instR191 (zll_main_multiply1785_inR47[128:1], zll_main_multiply1785_inR47[0], zll_main_multiply1785_outR47);
  assign zll_main_multiply1103_in = {zll_main_multiply1238_in[255:128], zll_main_multiply1238_in[127:0], zll_main_multiply1785_outR47};
  assign id_inR144 = zll_main_multiply1103_in[383:256];
  assign zll_main_multiply413_in = {zll_main_multiply1103_in[383:256], zll_main_multiply1103_in[255:128], zll_main_multiply1103_in[127:0], id_inR144[79]};
  assign id_inR145 = zll_main_multiply413_in[384:257];
  assign zll_main_multiply1792_inR48 = {zll_main_multiply413_in[256:129], id_inR145[79]};
  ZLL_Main_multiply1792  instR192 (zll_main_multiply1792_inR48[128:1], zll_main_multiply1792_inR48[0], zll_main_multiply1792_outR48);
  assign zll_main_multiply1749_inR22 = {zll_main_multiply413_in[256:129], zll_main_multiply413_in[128:1], zll_main_multiply413_in[0]};
  ZLL_Main_multiply1749  instR193 (zll_main_multiply1749_inR22[256:129], zll_main_multiply1749_inR22[128:1], zll_main_multiply1749_outR22);
  assign zll_main_multiply1177_in = {zll_main_multiply1103_in[383:256], zll_main_multiply1103_in[127:0], (zll_main_multiply1749_inR22[0] == 1'h1) ? zll_main_multiply1749_outR22 : zll_main_multiply1792_outR48};
  assign id_inR146 = zll_main_multiply1177_in[255:128];
  assign rewire_prelude_not_inR48 = id_inR146[0];
  ReWire_Prelude_not  instR194 (rewire_prelude_not_inR48[0], rewire_prelude_not_outR48);
  assign zll_main_multiply1785_inR48 = {zll_main_multiply1177_in[255:128], rewire_prelude_not_outR48};
  ZLL_Main_multiply1785  instR195 (zll_main_multiply1785_inR48[128:1], zll_main_multiply1785_inR48[0], zll_main_multiply1785_outR48);
  assign zll_main_multiply716_in = {zll_main_multiply1177_in[127:0], zll_main_multiply1177_in[383:256], zll_main_multiply1785_outR48};
  assign id_inR147 = zll_main_multiply716_in[255:128];
  assign zll_main_multiply384_in = {zll_main_multiply716_in[383:256], zll_main_multiply716_in[255:128], zll_main_multiply716_in[127:0], id_inR147[78]};
  assign id_inR148 = zll_main_multiply384_in[256:129];
  assign zll_main_multiply1792_inR49 = {zll_main_multiply384_in[384:257], id_inR148[78]};
  ZLL_Main_multiply1792  instR196 (zll_main_multiply1792_inR49[128:1], zll_main_multiply1792_inR49[0], zll_main_multiply1792_outR49);
  assign zll_main_multiply1749_inR23 = {zll_main_multiply384_in[384:257], zll_main_multiply384_in[128:1], zll_main_multiply384_in[0]};
  ZLL_Main_multiply1749  instR197 (zll_main_multiply1749_inR23[256:129], zll_main_multiply1749_inR23[128:1], zll_main_multiply1749_outR23);
  assign zll_main_multiply267_in = {zll_main_multiply716_in[255:128], zll_main_multiply716_in[127:0], (zll_main_multiply1749_inR23[0] == 1'h1) ? zll_main_multiply1749_outR23 : zll_main_multiply1792_outR49};
  assign id_inR149 = zll_main_multiply267_in[255:128];
  assign rewire_prelude_not_inR49 = id_inR149[0];
  ReWire_Prelude_not  instR198 (rewire_prelude_not_inR49[0], rewire_prelude_not_outR49);
  assign zll_main_multiply1785_inR49 = {zll_main_multiply267_in[255:128], rewire_prelude_not_outR49};
  ZLL_Main_multiply1785  instR199 (zll_main_multiply1785_inR49[128:1], zll_main_multiply1785_inR49[0], zll_main_multiply1785_outR49);
  assign zll_main_multiply72_in = {zll_main_multiply267_in[383:256], zll_main_multiply267_in[127:0], zll_main_multiply1785_outR49};
  assign id_inR150 = zll_main_multiply72_in[383:256];
  assign zll_main_multiply928_in = {zll_main_multiply72_in[127:0], zll_main_multiply72_in[383:256], zll_main_multiply72_in[255:128], id_inR150[77]};
  assign id_inR151 = zll_main_multiply928_in[256:129];
  assign zll_main_multiply1792_inR50 = {zll_main_multiply928_in[128:1], id_inR151[77]};
  ZLL_Main_multiply1792  instR200 (zll_main_multiply1792_inR50[128:1], zll_main_multiply1792_inR50[0], zll_main_multiply1792_outR50);
  assign zll_main_multiply1788_inR26 = {zll_main_multiply928_in[384:257], zll_main_multiply928_in[128:1], zll_main_multiply928_in[0]};
  ZLL_Main_multiply1788  instR201 (zll_main_multiply1788_inR26[256:129], zll_main_multiply1788_inR26[128:1], zll_main_multiply1788_outR26);
  assign zll_main_multiply849_in = {zll_main_multiply72_in[127:0], zll_main_multiply72_in[383:256], (zll_main_multiply1788_inR26[0] == 1'h1) ? zll_main_multiply1788_outR26 : zll_main_multiply1792_outR50};
  assign id_inR152 = zll_main_multiply849_in[383:256];
  assign rewire_prelude_not_inR50 = id_inR152[0];
  ReWire_Prelude_not  instR202 (rewire_prelude_not_inR50[0], rewire_prelude_not_outR50);
  assign zll_main_multiply1785_inR50 = {zll_main_multiply849_in[383:256], rewire_prelude_not_outR50};
  ZLL_Main_multiply1785  instR203 (zll_main_multiply1785_inR50[128:1], zll_main_multiply1785_inR50[0], zll_main_multiply1785_outR50);
  assign zll_main_multiply1488_in = {zll_main_multiply849_in[127:0], zll_main_multiply849_in[255:128], zll_main_multiply1785_outR50};
  assign id_inR153 = zll_main_multiply1488_in[255:128];
  assign zll_main_multiply996_in = {zll_main_multiply1488_in[383:256], zll_main_multiply1488_in[255:128], zll_main_multiply1488_in[127:0], id_inR153[76]};
  assign id_inR154 = zll_main_multiply996_in[256:129];
  assign zll_main_multiply1792_inR51 = {zll_main_multiply996_in[384:257], id_inR154[76]};
  ZLL_Main_multiply1792  instR204 (zll_main_multiply1792_inR51[128:1], zll_main_multiply1792_inR51[0], zll_main_multiply1792_outR51);
  assign zll_main_multiply1749_inR24 = {zll_main_multiply996_in[384:257], zll_main_multiply996_in[128:1], zll_main_multiply996_in[0]};
  ZLL_Main_multiply1749  instR205 (zll_main_multiply1749_inR24[256:129], zll_main_multiply1749_inR24[128:1], zll_main_multiply1749_outR24);
  assign zll_main_multiply287_in = {zll_main_multiply1488_in[255:128], zll_main_multiply1488_in[127:0], (zll_main_multiply1749_inR24[0] == 1'h1) ? zll_main_multiply1749_outR24 : zll_main_multiply1792_outR51};
  assign id_inR155 = zll_main_multiply287_in[255:128];
  assign rewire_prelude_not_inR51 = id_inR155[0];
  ReWire_Prelude_not  instR206 (rewire_prelude_not_inR51[0], rewire_prelude_not_outR51);
  assign zll_main_multiply1785_inR51 = {zll_main_multiply287_in[255:128], rewire_prelude_not_outR51};
  ZLL_Main_multiply1785  instR207 (zll_main_multiply1785_inR51[128:1], zll_main_multiply1785_inR51[0], zll_main_multiply1785_outR51);
  assign zll_main_multiply1648_in = {zll_main_multiply287_in[383:256], zll_main_multiply287_in[127:0], zll_main_multiply1785_outR51};
  assign id_inR156 = zll_main_multiply1648_in[383:256];
  assign zll_main_multiply868_in = {zll_main_multiply1648_in[383:256], zll_main_multiply1648_in[255:128], zll_main_multiply1648_in[127:0], id_inR156[75]};
  assign id_inR157 = zll_main_multiply868_in[384:257];
  assign zll_main_multiply1792_inR52 = {zll_main_multiply868_in[256:129], id_inR157[75]};
  ZLL_Main_multiply1792  instR208 (zll_main_multiply1792_inR52[128:1], zll_main_multiply1792_inR52[0], zll_main_multiply1792_outR52);
  assign zll_main_multiply1749_inR25 = {zll_main_multiply868_in[256:129], zll_main_multiply868_in[128:1], zll_main_multiply868_in[0]};
  ZLL_Main_multiply1749  instR209 (zll_main_multiply1749_inR25[256:129], zll_main_multiply1749_inR25[128:1], zll_main_multiply1749_outR25);
  assign zll_main_multiply594_in = {zll_main_multiply1648_in[383:256], zll_main_multiply1648_in[127:0], (zll_main_multiply1749_inR25[0] == 1'h1) ? zll_main_multiply1749_outR25 : zll_main_multiply1792_outR52};
  assign id_inR158 = zll_main_multiply594_in[255:128];
  assign rewire_prelude_not_inR52 = id_inR158[0];
  ReWire_Prelude_not  instR210 (rewire_prelude_not_inR52[0], rewire_prelude_not_outR52);
  assign zll_main_multiply1785_inR52 = {zll_main_multiply594_in[255:128], rewire_prelude_not_outR52};
  ZLL_Main_multiply1785  instR211 (zll_main_multiply1785_inR52[128:1], zll_main_multiply1785_inR52[0], zll_main_multiply1785_outR52);
  assign zll_main_multiply1745_in = {zll_main_multiply594_in[383:256], zll_main_multiply594_in[127:0], zll_main_multiply1785_outR52};
  assign id_inR159 = zll_main_multiply1745_in[383:256];
  assign zll_main_multiply976_in = {zll_main_multiply1745_in[127:0], zll_main_multiply1745_in[383:256], zll_main_multiply1745_in[255:128], id_inR159[74]};
  assign id_inR160 = zll_main_multiply976_in[256:129];
  assign zll_main_multiply1792_inR53 = {zll_main_multiply976_in[128:1], id_inR160[74]};
  ZLL_Main_multiply1792  instR212 (zll_main_multiply1792_inR53[128:1], zll_main_multiply1792_inR53[0], zll_main_multiply1792_outR53);
  assign zll_main_multiply1788_inR27 = {zll_main_multiply976_in[384:257], zll_main_multiply976_in[128:1], zll_main_multiply976_in[0]};
  ZLL_Main_multiply1788  instR213 (zll_main_multiply1788_inR27[256:129], zll_main_multiply1788_inR27[128:1], zll_main_multiply1788_outR27);
  assign zll_main_multiply436_in = {zll_main_multiply1745_in[127:0], zll_main_multiply1745_in[383:256], (zll_main_multiply1788_inR27[0] == 1'h1) ? zll_main_multiply1788_outR27 : zll_main_multiply1792_outR53};
  assign id_inR161 = zll_main_multiply436_in[383:256];
  assign rewire_prelude_not_inR53 = id_inR161[0];
  ReWire_Prelude_not  instR214 (rewire_prelude_not_inR53[0], rewire_prelude_not_outR53);
  assign zll_main_multiply1785_inR53 = {zll_main_multiply436_in[383:256], rewire_prelude_not_outR53};
  ZLL_Main_multiply1785  instR215 (zll_main_multiply1785_inR53[128:1], zll_main_multiply1785_inR53[0], zll_main_multiply1785_outR53);
  assign zll_main_multiply260_in = {zll_main_multiply436_in[255:128], zll_main_multiply436_in[127:0], zll_main_multiply1785_outR53};
  assign id_inR162 = zll_main_multiply260_in[383:256];
  assign zll_main_multiply1381_in = {zll_main_multiply260_in[383:256], zll_main_multiply260_in[127:0], zll_main_multiply260_in[255:128], id_inR162[73]};
  assign id_inR163 = zll_main_multiply1381_in[384:257];
  assign zll_main_multiply1792_inR54 = {zll_main_multiply1381_in[128:1], id_inR163[73]};
  ZLL_Main_multiply1792  instR216 (zll_main_multiply1792_inR54[128:1], zll_main_multiply1792_inR54[0], zll_main_multiply1792_outR54);
  assign zll_main_multiply1788_inR28 = {zll_main_multiply1381_in[256:129], zll_main_multiply1381_in[128:1], zll_main_multiply1381_in[0]};
  ZLL_Main_multiply1788  instR217 (zll_main_multiply1788_inR28[256:129], zll_main_multiply1788_inR28[128:1], zll_main_multiply1788_outR28);
  assign zll_main_multiply1598_in = {zll_main_multiply260_in[383:256], zll_main_multiply260_in[127:0], (zll_main_multiply1788_inR28[0] == 1'h1) ? zll_main_multiply1788_outR28 : zll_main_multiply1792_outR54};
  assign id_inR164 = zll_main_multiply1598_in[255:128];
  assign rewire_prelude_not_inR54 = id_inR164[0];
  ReWire_Prelude_not  instR218 (rewire_prelude_not_inR54[0], rewire_prelude_not_outR54);
  assign zll_main_multiply1785_inR54 = {zll_main_multiply1598_in[255:128], rewire_prelude_not_outR54};
  ZLL_Main_multiply1785  instR219 (zll_main_multiply1785_inR54[128:1], zll_main_multiply1785_inR54[0], zll_main_multiply1785_outR54);
  assign zll_main_multiply1610_in = {zll_main_multiply1598_in[383:256], zll_main_multiply1598_in[127:0], zll_main_multiply1785_outR54};
  assign id_inR165 = zll_main_multiply1610_in[383:256];
  assign zll_main_multiply806_in = {zll_main_multiply1610_in[127:0], zll_main_multiply1610_in[383:256], zll_main_multiply1610_in[255:128], id_inR165[72]};
  assign id_inR166 = zll_main_multiply806_in[256:129];
  assign zll_main_multiply1792_inR55 = {zll_main_multiply806_in[128:1], id_inR166[72]};
  ZLL_Main_multiply1792  instR220 (zll_main_multiply1792_inR55[128:1], zll_main_multiply1792_inR55[0], zll_main_multiply1792_outR55);
  assign zll_main_multiply1788_inR29 = {zll_main_multiply806_in[384:257], zll_main_multiply806_in[128:1], zll_main_multiply806_in[0]};
  ZLL_Main_multiply1788  instR221 (zll_main_multiply1788_inR29[256:129], zll_main_multiply1788_inR29[128:1], zll_main_multiply1788_outR29);
  assign zll_main_multiply830_in = {zll_main_multiply1610_in[127:0], zll_main_multiply1610_in[383:256], (zll_main_multiply1788_inR29[0] == 1'h1) ? zll_main_multiply1788_outR29 : zll_main_multiply1792_outR55};
  assign id_inR167 = zll_main_multiply830_in[383:256];
  assign rewire_prelude_not_inR55 = id_inR167[0];
  ReWire_Prelude_not  instR222 (rewire_prelude_not_inR55[0], rewire_prelude_not_outR55);
  assign zll_main_multiply1785_inR55 = {zll_main_multiply830_in[383:256], rewire_prelude_not_outR55};
  ZLL_Main_multiply1785  instR223 (zll_main_multiply1785_inR55[128:1], zll_main_multiply1785_inR55[0], zll_main_multiply1785_outR55);
  assign zll_main_multiply792_in = {zll_main_multiply830_in[127:0], zll_main_multiply830_in[255:128], zll_main_multiply1785_outR55};
  assign id_inR168 = zll_main_multiply792_in[255:128];
  assign zll_main_multiply1584_in = {zll_main_multiply792_in[383:256], zll_main_multiply792_in[255:128], zll_main_multiply792_in[127:0], id_inR168[71]};
  assign id_inR169 = zll_main_multiply1584_in[256:129];
  assign zll_main_multiply1792_inR56 = {zll_main_multiply1584_in[384:257], id_inR169[71]};
  ZLL_Main_multiply1792  instR224 (zll_main_multiply1792_inR56[128:1], zll_main_multiply1792_inR56[0], zll_main_multiply1792_outR56);
  assign zll_main_multiply1749_inR26 = {zll_main_multiply1584_in[384:257], zll_main_multiply1584_in[128:1], zll_main_multiply1584_in[0]};
  ZLL_Main_multiply1749  instR225 (zll_main_multiply1749_inR26[256:129], zll_main_multiply1749_inR26[128:1], zll_main_multiply1749_outR26);
  assign zll_main_multiply14_in = {zll_main_multiply792_in[255:128], zll_main_multiply792_in[127:0], (zll_main_multiply1749_inR26[0] == 1'h1) ? zll_main_multiply1749_outR26 : zll_main_multiply1792_outR56};
  assign id_inR170 = zll_main_multiply14_in[255:128];
  assign rewire_prelude_not_inR56 = id_inR170[0];
  ReWire_Prelude_not  instR226 (rewire_prelude_not_inR56[0], rewire_prelude_not_outR56);
  assign zll_main_multiply1785_inR56 = {zll_main_multiply14_in[255:128], rewire_prelude_not_outR56};
  ZLL_Main_multiply1785  instR227 (zll_main_multiply1785_inR56[128:1], zll_main_multiply1785_inR56[0], zll_main_multiply1785_outR56);
  assign zll_main_multiply1099_in = {zll_main_multiply14_in[127:0], zll_main_multiply14_in[383:256], zll_main_multiply1785_outR56};
  assign id_inR171 = zll_main_multiply1099_in[255:128];
  assign zll_main_multiply719_in = {zll_main_multiply1099_in[383:256], zll_main_multiply1099_in[255:128], zll_main_multiply1099_in[127:0], id_inR171[70]};
  assign id_inR172 = zll_main_multiply719_in[256:129];
  assign zll_main_multiply1792_inR57 = {zll_main_multiply719_in[384:257], id_inR172[70]};
  ZLL_Main_multiply1792  instR228 (zll_main_multiply1792_inR57[128:1], zll_main_multiply1792_inR57[0], zll_main_multiply1792_outR57);
  assign zll_main_multiply1749_inR27 = {zll_main_multiply719_in[384:257], zll_main_multiply719_in[128:1], zll_main_multiply719_in[0]};
  ZLL_Main_multiply1749  instR229 (zll_main_multiply1749_inR27[256:129], zll_main_multiply1749_inR27[128:1], zll_main_multiply1749_outR27);
  assign zll_main_multiply150_in = {zll_main_multiply1099_in[255:128], zll_main_multiply1099_in[127:0], (zll_main_multiply1749_inR27[0] == 1'h1) ? zll_main_multiply1749_outR27 : zll_main_multiply1792_outR57};
  assign id_inR173 = zll_main_multiply150_in[255:128];
  assign rewire_prelude_not_inR57 = id_inR173[0];
  ReWire_Prelude_not  instR230 (rewire_prelude_not_inR57[0], rewire_prelude_not_outR57);
  assign zll_main_multiply1785_inR57 = {zll_main_multiply150_in[255:128], rewire_prelude_not_outR57};
  ZLL_Main_multiply1785  instR231 (zll_main_multiply1785_inR57[128:1], zll_main_multiply1785_inR57[0], zll_main_multiply1785_outR57);
  assign zll_main_multiply1791_in = {zll_main_multiply150_in[383:256], zll_main_multiply150_in[127:0], zll_main_multiply1785_outR57};
  assign id_inR174 = zll_main_multiply1791_in[383:256];
  assign zll_main_multiply472_in = {zll_main_multiply1791_in[383:256], zll_main_multiply1791_in[255:128], zll_main_multiply1791_in[127:0], id_inR174[69]};
  assign id_inR175 = zll_main_multiply472_in[384:257];
  assign zll_main_multiply1792_inR58 = {zll_main_multiply472_in[256:129], id_inR175[69]};
  ZLL_Main_multiply1792  instR232 (zll_main_multiply1792_inR58[128:1], zll_main_multiply1792_inR58[0], zll_main_multiply1792_outR58);
  assign zll_main_multiply1749_inR28 = {zll_main_multiply472_in[256:129], zll_main_multiply472_in[128:1], zll_main_multiply472_in[0]};
  ZLL_Main_multiply1749  instR233 (zll_main_multiply1749_inR28[256:129], zll_main_multiply1749_inR28[128:1], zll_main_multiply1749_outR28);
  assign zll_main_multiply1270_in = {zll_main_multiply1791_in[383:256], zll_main_multiply1791_in[127:0], (zll_main_multiply1749_inR28[0] == 1'h1) ? zll_main_multiply1749_outR28 : zll_main_multiply1792_outR58};
  assign id_inR176 = zll_main_multiply1270_in[255:128];
  assign rewire_prelude_not_inR58 = id_inR176[0];
  ReWire_Prelude_not  instR234 (rewire_prelude_not_inR58[0], rewire_prelude_not_outR58);
  assign zll_main_multiply1785_inR58 = {zll_main_multiply1270_in[255:128], rewire_prelude_not_outR58};
  ZLL_Main_multiply1785  instR235 (zll_main_multiply1785_inR58[128:1], zll_main_multiply1785_inR58[0], zll_main_multiply1785_outR58);
  assign zll_main_multiply1207_in = {zll_main_multiply1270_in[383:256], zll_main_multiply1270_in[127:0], zll_main_multiply1785_outR58};
  assign id_inR177 = zll_main_multiply1207_in[383:256];
  assign zll_main_multiply1210_in = {zll_main_multiply1207_in[127:0], zll_main_multiply1207_in[383:256], zll_main_multiply1207_in[255:128], id_inR177[68]};
  assign id_inR178 = zll_main_multiply1210_in[256:129];
  assign zll_main_multiply1792_inR59 = {zll_main_multiply1210_in[128:1], id_inR178[68]};
  ZLL_Main_multiply1792  instR236 (zll_main_multiply1792_inR59[128:1], zll_main_multiply1792_inR59[0], zll_main_multiply1792_outR59);
  assign zll_main_multiply1788_inR30 = {zll_main_multiply1210_in[384:257], zll_main_multiply1210_in[128:1], zll_main_multiply1210_in[0]};
  ZLL_Main_multiply1788  instR237 (zll_main_multiply1788_inR30[256:129], zll_main_multiply1788_inR30[128:1], zll_main_multiply1788_outR30);
  assign zll_main_multiply215_in = {zll_main_multiply1207_in[127:0], zll_main_multiply1207_in[383:256], (zll_main_multiply1788_inR30[0] == 1'h1) ? zll_main_multiply1788_outR30 : zll_main_multiply1792_outR59};
  assign id_inR179 = zll_main_multiply215_in[383:256];
  assign rewire_prelude_not_inR59 = id_inR179[0];
  ReWire_Prelude_not  instR238 (rewire_prelude_not_inR59[0], rewire_prelude_not_outR59);
  assign zll_main_multiply1785_inR59 = {zll_main_multiply215_in[383:256], rewire_prelude_not_outR59};
  ZLL_Main_multiply1785  instR239 (zll_main_multiply1785_inR59[128:1], zll_main_multiply1785_inR59[0], zll_main_multiply1785_outR59);
  assign zll_main_multiply1202_in = {zll_main_multiply215_in[255:128], zll_main_multiply215_in[127:0], zll_main_multiply1785_outR59};
  assign id_inR180 = zll_main_multiply1202_in[383:256];
  assign zll_main_multiply28_in = {zll_main_multiply1202_in[383:256], zll_main_multiply1202_in[255:128], zll_main_multiply1202_in[127:0], id_inR180[67]};
  assign id_inR181 = zll_main_multiply28_in[384:257];
  assign zll_main_multiply1792_inR60 = {zll_main_multiply28_in[256:129], id_inR181[67]};
  ZLL_Main_multiply1792  instR240 (zll_main_multiply1792_inR60[128:1], zll_main_multiply1792_inR60[0], zll_main_multiply1792_outR60);
  assign zll_main_multiply1749_inR29 = {zll_main_multiply28_in[256:129], zll_main_multiply28_in[128:1], zll_main_multiply28_in[0]};
  ZLL_Main_multiply1749  instR241 (zll_main_multiply1749_inR29[256:129], zll_main_multiply1749_inR29[128:1], zll_main_multiply1749_outR29);
  assign zll_main_multiply9_in = {zll_main_multiply1202_in[383:256], zll_main_multiply1202_in[127:0], (zll_main_multiply1749_inR29[0] == 1'h1) ? zll_main_multiply1749_outR29 : zll_main_multiply1792_outR60};
  assign id_inR182 = zll_main_multiply9_in[255:128];
  assign rewire_prelude_not_inR60 = id_inR182[0];
  ReWire_Prelude_not  instR242 (rewire_prelude_not_inR60[0], rewire_prelude_not_outR60);
  assign zll_main_multiply1785_inR60 = {zll_main_multiply9_in[255:128], rewire_prelude_not_outR60};
  ZLL_Main_multiply1785  instR243 (zll_main_multiply1785_inR60[128:1], zll_main_multiply1785_inR60[0], zll_main_multiply1785_outR60);
  assign zll_main_multiply1279_in = {zll_main_multiply9_in[127:0], zll_main_multiply9_in[383:256], zll_main_multiply1785_outR60};
  assign id_inR183 = zll_main_multiply1279_in[255:128];
  assign zll_main_multiply132_in = {zll_main_multiply1279_in[383:256], zll_main_multiply1279_in[255:128], zll_main_multiply1279_in[127:0], id_inR183[66]};
  assign id_inR184 = zll_main_multiply132_in[256:129];
  assign zll_main_multiply1792_inR61 = {zll_main_multiply132_in[384:257], id_inR184[66]};
  ZLL_Main_multiply1792  instR244 (zll_main_multiply1792_inR61[128:1], zll_main_multiply1792_inR61[0], zll_main_multiply1792_outR61);
  assign zll_main_multiply1749_inR30 = {zll_main_multiply132_in[384:257], zll_main_multiply132_in[128:1], zll_main_multiply132_in[0]};
  ZLL_Main_multiply1749  instR245 (zll_main_multiply1749_inR30[256:129], zll_main_multiply1749_inR30[128:1], zll_main_multiply1749_outR30);
  assign zll_main_multiply530_in = {zll_main_multiply1279_in[255:128], zll_main_multiply1279_in[127:0], (zll_main_multiply1749_inR30[0] == 1'h1) ? zll_main_multiply1749_outR30 : zll_main_multiply1792_outR61};
  assign id_inR185 = zll_main_multiply530_in[255:128];
  assign rewire_prelude_not_inR61 = id_inR185[0];
  ReWire_Prelude_not  instR246 (rewire_prelude_not_inR61[0], rewire_prelude_not_outR61);
  assign zll_main_multiply1785_inR61 = {zll_main_multiply530_in[255:128], rewire_prelude_not_outR61};
  ZLL_Main_multiply1785  instR247 (zll_main_multiply1785_inR61[128:1], zll_main_multiply1785_inR61[0], zll_main_multiply1785_outR61);
  assign zll_main_multiply1445_in = {zll_main_multiply530_in[127:0], zll_main_multiply530_in[383:256], zll_main_multiply1785_outR61};
  assign id_inR186 = zll_main_multiply1445_in[255:128];
  assign zll_main_multiply1545_in = {zll_main_multiply1445_in[127:0], zll_main_multiply1445_in[383:256], zll_main_multiply1445_in[255:128], id_inR186[65]};
  assign id_inR187 = zll_main_multiply1545_in[128:1];
  assign zll_main_multiply1792_inR62 = {zll_main_multiply1545_in[256:129], id_inR187[65]};
  ZLL_Main_multiply1792  instR248 (zll_main_multiply1792_inR62[128:1], zll_main_multiply1792_inR62[0], zll_main_multiply1792_outR62);
  assign zll_main_multiply1788_inR31 = {zll_main_multiply1545_in[384:257], zll_main_multiply1545_in[256:129], zll_main_multiply1545_in[0]};
  ZLL_Main_multiply1788  instR249 (zll_main_multiply1788_inR31[256:129], zll_main_multiply1788_inR31[128:1], zll_main_multiply1788_outR31);
  assign zll_main_multiply1517_in = {zll_main_multiply1445_in[127:0], zll_main_multiply1445_in[255:128], (zll_main_multiply1788_inR31[0] == 1'h1) ? zll_main_multiply1788_outR31 : zll_main_multiply1792_outR62};
  assign id_inR188 = zll_main_multiply1517_in[383:256];
  assign rewire_prelude_not_inR62 = id_inR188[0];
  ReWire_Prelude_not  instR250 (rewire_prelude_not_inR62[0], rewire_prelude_not_outR62);
  assign zll_main_multiply1785_inR62 = {zll_main_multiply1517_in[383:256], rewire_prelude_not_outR62};
  ZLL_Main_multiply1785  instR251 (zll_main_multiply1785_inR62[128:1], zll_main_multiply1785_inR62[0], zll_main_multiply1785_outR62);
  assign zll_main_multiply326_in = {zll_main_multiply1517_in[255:128], zll_main_multiply1517_in[127:0], zll_main_multiply1785_outR62};
  assign id_inR189 = zll_main_multiply326_in[383:256];
  assign zll_main_multiply1468_in = {zll_main_multiply326_in[127:0], zll_main_multiply326_in[383:256], zll_main_multiply326_in[255:128], id_inR189[64]};
  assign id_inR190 = zll_main_multiply1468_in[256:129];
  assign zll_main_multiply1792_inR63 = {zll_main_multiply1468_in[128:1], id_inR190[64]};
  ZLL_Main_multiply1792  instR252 (zll_main_multiply1792_inR63[128:1], zll_main_multiply1792_inR63[0], zll_main_multiply1792_outR63);
  assign zll_main_multiply1788_inR32 = {zll_main_multiply1468_in[384:257], zll_main_multiply1468_in[128:1], zll_main_multiply1468_in[0]};
  ZLL_Main_multiply1788  instR253 (zll_main_multiply1788_inR32[256:129], zll_main_multiply1788_inR32[128:1], zll_main_multiply1788_outR32);
  assign zll_main_multiply1693_in = {zll_main_multiply326_in[127:0], zll_main_multiply326_in[383:256], (zll_main_multiply1788_inR32[0] == 1'h1) ? zll_main_multiply1788_outR32 : zll_main_multiply1792_outR63};
  assign id_inR191 = zll_main_multiply1693_in[383:256];
  assign rewire_prelude_not_inR63 = id_inR191[0];
  ReWire_Prelude_not  instR254 (rewire_prelude_not_inR63[0], rewire_prelude_not_outR63);
  assign zll_main_multiply1785_inR63 = {zll_main_multiply1693_in[383:256], rewire_prelude_not_outR63};
  ZLL_Main_multiply1785  instR255 (zll_main_multiply1785_inR63[128:1], zll_main_multiply1785_inR63[0], zll_main_multiply1785_outR63);
  assign zll_main_multiply284_in = {zll_main_multiply1693_in[255:128], zll_main_multiply1693_in[127:0], zll_main_multiply1785_outR63};
  assign id_inR192 = zll_main_multiply284_in[383:256];
  assign zll_main_multiply1639_in = {zll_main_multiply284_in[127:0], zll_main_multiply284_in[383:256], zll_main_multiply284_in[255:128], id_inR192[63]};
  assign id_inR193 = zll_main_multiply1639_in[256:129];
  assign zll_main_multiply1792_inR64 = {zll_main_multiply1639_in[128:1], id_inR193[63]};
  ZLL_Main_multiply1792  instR256 (zll_main_multiply1792_inR64[128:1], zll_main_multiply1792_inR64[0], zll_main_multiply1792_outR64);
  assign zll_main_multiply1788_inR33 = {zll_main_multiply1639_in[384:257], zll_main_multiply1639_in[128:1], zll_main_multiply1639_in[0]};
  ZLL_Main_multiply1788  instR257 (zll_main_multiply1788_inR33[256:129], zll_main_multiply1788_inR33[128:1], zll_main_multiply1788_outR33);
  assign zll_main_multiply675_in = {zll_main_multiply284_in[127:0], zll_main_multiply284_in[383:256], (zll_main_multiply1788_inR33[0] == 1'h1) ? zll_main_multiply1788_outR33 : zll_main_multiply1792_outR64};
  assign id_inR194 = zll_main_multiply675_in[383:256];
  assign rewire_prelude_not_inR64 = id_inR194[0];
  ReWire_Prelude_not  instR258 (rewire_prelude_not_inR64[0], rewire_prelude_not_outR64);
  assign zll_main_multiply1785_inR64 = {zll_main_multiply675_in[383:256], rewire_prelude_not_outR64};
  ZLL_Main_multiply1785  instR259 (zll_main_multiply1785_inR64[128:1], zll_main_multiply1785_inR64[0], zll_main_multiply1785_outR64);
  assign zll_main_multiply1633_in = {zll_main_multiply675_in[127:0], zll_main_multiply675_in[255:128], zll_main_multiply1785_outR64};
  assign id_inR195 = zll_main_multiply1633_in[255:128];
  assign zll_main_multiply1469_in = {zll_main_multiply1633_in[383:256], zll_main_multiply1633_in[255:128], zll_main_multiply1633_in[127:0], id_inR195[62]};
  assign id_inR196 = zll_main_multiply1469_in[256:129];
  assign zll_main_multiply1792_inR65 = {zll_main_multiply1469_in[384:257], id_inR196[62]};
  ZLL_Main_multiply1792  instR260 (zll_main_multiply1792_inR65[128:1], zll_main_multiply1792_inR65[0], zll_main_multiply1792_outR65);
  assign zll_main_multiply1749_inR31 = {zll_main_multiply1469_in[384:257], zll_main_multiply1469_in[128:1], zll_main_multiply1469_in[0]};
  ZLL_Main_multiply1749  instR261 (zll_main_multiply1749_inR31[256:129], zll_main_multiply1749_inR31[128:1], zll_main_multiply1749_outR31);
  assign zll_main_multiply300_in = {zll_main_multiply1633_in[255:128], zll_main_multiply1633_in[127:0], (zll_main_multiply1749_inR31[0] == 1'h1) ? zll_main_multiply1749_outR31 : zll_main_multiply1792_outR65};
  assign id_inR197 = zll_main_multiply300_in[255:128];
  assign rewire_prelude_not_inR65 = id_inR197[0];
  ReWire_Prelude_not  instR262 (rewire_prelude_not_inR65[0], rewire_prelude_not_outR65);
  assign zll_main_multiply1785_inR65 = {zll_main_multiply300_in[255:128], rewire_prelude_not_outR65};
  ZLL_Main_multiply1785  instR263 (zll_main_multiply1785_inR65[128:1], zll_main_multiply1785_inR65[0], zll_main_multiply1785_outR65);
  assign zll_main_multiply1709_in = {zll_main_multiply300_in[127:0], zll_main_multiply300_in[383:256], zll_main_multiply1785_outR65};
  assign id_inR198 = zll_main_multiply1709_in[255:128];
  assign zll_main_multiply1_in = {zll_main_multiply1709_in[127:0], zll_main_multiply1709_in[383:256], zll_main_multiply1709_in[255:128], id_inR198[61]};
  assign id_inR199 = zll_main_multiply1_in[128:1];
  assign zll_main_multiply1792_inR66 = {zll_main_multiply1_in[256:129], id_inR199[61]};
  ZLL_Main_multiply1792  instR264 (zll_main_multiply1792_inR66[128:1], zll_main_multiply1792_inR66[0], zll_main_multiply1792_outR66);
  assign zll_main_multiply1788_inR34 = {zll_main_multiply1_in[384:257], zll_main_multiply1_in[256:129], zll_main_multiply1_in[0]};
  ZLL_Main_multiply1788  instR265 (zll_main_multiply1788_inR34[256:129], zll_main_multiply1788_inR34[128:1], zll_main_multiply1788_outR34);
  assign zll_main_multiply837_in = {zll_main_multiply1709_in[127:0], zll_main_multiply1709_in[255:128], (zll_main_multiply1788_inR34[0] == 1'h1) ? zll_main_multiply1788_outR34 : zll_main_multiply1792_outR66};
  assign id_inR200 = zll_main_multiply837_in[383:256];
  assign rewire_prelude_not_inR66 = id_inR200[0];
  ReWire_Prelude_not  instR266 (rewire_prelude_not_inR66[0], rewire_prelude_not_outR66);
  assign zll_main_multiply1785_inR66 = {zll_main_multiply837_in[383:256], rewire_prelude_not_outR66};
  ZLL_Main_multiply1785  instR267 (zll_main_multiply1785_inR66[128:1], zll_main_multiply1785_inR66[0], zll_main_multiply1785_outR66);
  assign zll_main_multiply714_in = {zll_main_multiply837_in[127:0], zll_main_multiply837_in[255:128], zll_main_multiply1785_outR66};
  assign id_inR201 = zll_main_multiply714_in[255:128];
  assign zll_main_multiply1098_in = {zll_main_multiply714_in[383:256], zll_main_multiply714_in[255:128], zll_main_multiply714_in[127:0], id_inR201[60]};
  assign id_inR202 = zll_main_multiply1098_in[256:129];
  assign zll_main_multiply1792_inR67 = {zll_main_multiply1098_in[384:257], id_inR202[60]};
  ZLL_Main_multiply1792  instR268 (zll_main_multiply1792_inR67[128:1], zll_main_multiply1792_inR67[0], zll_main_multiply1792_outR67);
  assign zll_main_multiply1749_inR32 = {zll_main_multiply1098_in[384:257], zll_main_multiply1098_in[128:1], zll_main_multiply1098_in[0]};
  ZLL_Main_multiply1749  instR269 (zll_main_multiply1749_inR32[256:129], zll_main_multiply1749_inR32[128:1], zll_main_multiply1749_outR32);
  assign zll_main_multiply940_in = {zll_main_multiply714_in[255:128], zll_main_multiply714_in[127:0], (zll_main_multiply1749_inR32[0] == 1'h1) ? zll_main_multiply1749_outR32 : zll_main_multiply1792_outR67};
  assign id_inR203 = zll_main_multiply940_in[255:128];
  assign rewire_prelude_not_inR67 = id_inR203[0];
  ReWire_Prelude_not  instR270 (rewire_prelude_not_inR67[0], rewire_prelude_not_outR67);
  assign zll_main_multiply1785_inR67 = {zll_main_multiply940_in[255:128], rewire_prelude_not_outR67};
  ZLL_Main_multiply1785  instR271 (zll_main_multiply1785_inR67[128:1], zll_main_multiply1785_inR67[0], zll_main_multiply1785_outR67);
  assign zll_main_multiply76_in = {zll_main_multiply940_in[383:256], zll_main_multiply940_in[127:0], zll_main_multiply1785_outR67};
  assign id_inR204 = zll_main_multiply76_in[383:256];
  assign zll_main_multiply344_in = {zll_main_multiply76_in[127:0], zll_main_multiply76_in[383:256], zll_main_multiply76_in[255:128], id_inR204[59]};
  assign id_inR205 = zll_main_multiply344_in[256:129];
  assign zll_main_multiply1792_inR68 = {zll_main_multiply344_in[128:1], id_inR205[59]};
  ZLL_Main_multiply1792  instR272 (zll_main_multiply1792_inR68[128:1], zll_main_multiply1792_inR68[0], zll_main_multiply1792_outR68);
  assign zll_main_multiply1788_inR35 = {zll_main_multiply344_in[384:257], zll_main_multiply344_in[128:1], zll_main_multiply344_in[0]};
  ZLL_Main_multiply1788  instR273 (zll_main_multiply1788_inR35[256:129], zll_main_multiply1788_inR35[128:1], zll_main_multiply1788_outR35);
  assign zll_main_multiply970_in = {zll_main_multiply76_in[127:0], zll_main_multiply76_in[383:256], (zll_main_multiply1788_inR35[0] == 1'h1) ? zll_main_multiply1788_outR35 : zll_main_multiply1792_outR68};
  assign id_inR206 = zll_main_multiply970_in[383:256];
  assign rewire_prelude_not_inR68 = id_inR206[0];
  ReWire_Prelude_not  instR274 (rewire_prelude_not_inR68[0], rewire_prelude_not_outR68);
  assign zll_main_multiply1785_inR68 = {zll_main_multiply970_in[383:256], rewire_prelude_not_outR68};
  ZLL_Main_multiply1785  instR275 (zll_main_multiply1785_inR68[128:1], zll_main_multiply1785_inR68[0], zll_main_multiply1785_outR68);
  assign zll_main_multiply1765_in = {zll_main_multiply970_in[255:128], zll_main_multiply970_in[127:0], zll_main_multiply1785_outR68};
  assign id_inR207 = zll_main_multiply1765_in[383:256];
  assign zll_main_multiply1336_in = {zll_main_multiply1765_in[127:0], zll_main_multiply1765_in[383:256], zll_main_multiply1765_in[255:128], id_inR207[58]};
  assign id_inR208 = zll_main_multiply1336_in[256:129];
  assign zll_main_multiply1792_inR69 = {zll_main_multiply1336_in[128:1], id_inR208[58]};
  ZLL_Main_multiply1792  instR276 (zll_main_multiply1792_inR69[128:1], zll_main_multiply1792_inR69[0], zll_main_multiply1792_outR69);
  assign zll_main_multiply1788_inR36 = {zll_main_multiply1336_in[384:257], zll_main_multiply1336_in[128:1], zll_main_multiply1336_in[0]};
  ZLL_Main_multiply1788  instR277 (zll_main_multiply1788_inR36[256:129], zll_main_multiply1788_inR36[128:1], zll_main_multiply1788_outR36);
  assign zll_main_multiply1781_in = {zll_main_multiply1765_in[127:0], zll_main_multiply1765_in[383:256], (zll_main_multiply1788_inR36[0] == 1'h1) ? zll_main_multiply1788_outR36 : zll_main_multiply1792_outR69};
  assign id_inR209 = zll_main_multiply1781_in[383:256];
  assign rewire_prelude_not_inR69 = id_inR209[0];
  ReWire_Prelude_not  instR278 (rewire_prelude_not_inR69[0], rewire_prelude_not_outR69);
  assign zll_main_multiply1785_inR69 = {zll_main_multiply1781_in[383:256], rewire_prelude_not_outR69};
  ZLL_Main_multiply1785  instR279 (zll_main_multiply1785_inR69[128:1], zll_main_multiply1785_inR69[0], zll_main_multiply1785_outR69);
  assign zll_main_multiply1657_in = {zll_main_multiply1781_in[127:0], zll_main_multiply1781_in[255:128], zll_main_multiply1785_outR69};
  assign id_inR210 = zll_main_multiply1657_in[255:128];
  assign zll_main_multiply630_in = {zll_main_multiply1657_in[383:256], zll_main_multiply1657_in[255:128], zll_main_multiply1657_in[127:0], id_inR210[57]};
  assign id_inR211 = zll_main_multiply630_in[256:129];
  assign zll_main_multiply1792_inR70 = {zll_main_multiply630_in[384:257], id_inR211[57]};
  ZLL_Main_multiply1792  instR280 (zll_main_multiply1792_inR70[128:1], zll_main_multiply1792_inR70[0], zll_main_multiply1792_outR70);
  assign zll_main_multiply1749_inR33 = {zll_main_multiply630_in[384:257], zll_main_multiply630_in[128:1], zll_main_multiply630_in[0]};
  ZLL_Main_multiply1749  instR281 (zll_main_multiply1749_inR33[256:129], zll_main_multiply1749_inR33[128:1], zll_main_multiply1749_outR33);
  assign zll_main_multiply1717_in = {zll_main_multiply1657_in[255:128], zll_main_multiply1657_in[127:0], (zll_main_multiply1749_inR33[0] == 1'h1) ? zll_main_multiply1749_outR33 : zll_main_multiply1792_outR70};
  assign id_inR212 = zll_main_multiply1717_in[255:128];
  assign rewire_prelude_not_inR70 = id_inR212[0];
  ReWire_Prelude_not  instR282 (rewire_prelude_not_inR70[0], rewire_prelude_not_outR70);
  assign zll_main_multiply1785_inR70 = {zll_main_multiply1717_in[255:128], rewire_prelude_not_outR70};
  ZLL_Main_multiply1785  instR283 (zll_main_multiply1785_inR70[128:1], zll_main_multiply1785_inR70[0], zll_main_multiply1785_outR70);
  assign zll_main_multiply482_in = {zll_main_multiply1717_in[127:0], zll_main_multiply1717_in[383:256], zll_main_multiply1785_outR70};
  assign id_inR213 = zll_main_multiply482_in[255:128];
  assign zll_main_multiply1158_in = {zll_main_multiply482_in[127:0], zll_main_multiply482_in[383:256], zll_main_multiply482_in[255:128], id_inR213[56]};
  assign id_inR214 = zll_main_multiply1158_in[128:1];
  assign zll_main_multiply1792_inR71 = {zll_main_multiply1158_in[256:129], id_inR214[56]};
  ZLL_Main_multiply1792  instR284 (zll_main_multiply1792_inR71[128:1], zll_main_multiply1792_inR71[0], zll_main_multiply1792_outR71);
  assign zll_main_multiply1788_inR37 = {zll_main_multiply1158_in[384:257], zll_main_multiply1158_in[256:129], zll_main_multiply1158_in[0]};
  ZLL_Main_multiply1788  instR285 (zll_main_multiply1788_inR37[256:129], zll_main_multiply1788_inR37[128:1], zll_main_multiply1788_outR37);
  assign zll_main_multiply281_in = {zll_main_multiply482_in[127:0], zll_main_multiply482_in[255:128], (zll_main_multiply1788_inR37[0] == 1'h1) ? zll_main_multiply1788_outR37 : zll_main_multiply1792_outR71};
  assign id_inR215 = zll_main_multiply281_in[383:256];
  assign rewire_prelude_not_inR71 = id_inR215[0];
  ReWire_Prelude_not  instR286 (rewire_prelude_not_inR71[0], rewire_prelude_not_outR71);
  assign zll_main_multiply1785_inR71 = {zll_main_multiply281_in[383:256], rewire_prelude_not_outR71};
  ZLL_Main_multiply1785  instR287 (zll_main_multiply1785_inR71[128:1], zll_main_multiply1785_inR71[0], zll_main_multiply1785_outR71);
  assign zll_main_multiply1720_in = {zll_main_multiply281_in[127:0], zll_main_multiply281_in[255:128], zll_main_multiply1785_outR71};
  assign id_inR216 = zll_main_multiply1720_in[255:128];
  assign zll_main_multiply1640_in = {zll_main_multiply1720_in[383:256], zll_main_multiply1720_in[127:0], zll_main_multiply1720_in[255:128], id_inR216[55]};
  assign id_inR217 = zll_main_multiply1640_in[128:1];
  assign zll_main_multiply1792_inR72 = {zll_main_multiply1640_in[384:257], id_inR217[55]};
  ZLL_Main_multiply1792  instR288 (zll_main_multiply1792_inR72[128:1], zll_main_multiply1792_inR72[0], zll_main_multiply1792_outR72);
  assign zll_main_multiply1749_inR34 = {zll_main_multiply1640_in[384:257], zll_main_multiply1640_in[256:129], zll_main_multiply1640_in[0]};
  ZLL_Main_multiply1749  instR289 (zll_main_multiply1749_inR34[256:129], zll_main_multiply1749_inR34[128:1], zll_main_multiply1749_outR34);
  assign zll_main_multiply268_in = {zll_main_multiply1720_in[127:0], zll_main_multiply1720_in[255:128], (zll_main_multiply1749_inR34[0] == 1'h1) ? zll_main_multiply1749_outR34 : zll_main_multiply1792_outR72};
  assign id_inR218 = zll_main_multiply268_in[383:256];
  assign rewire_prelude_not_inR72 = id_inR218[0];
  ReWire_Prelude_not  instR290 (rewire_prelude_not_inR72[0], rewire_prelude_not_outR72);
  assign zll_main_multiply1785_inR72 = {zll_main_multiply268_in[383:256], rewire_prelude_not_outR72};
  ZLL_Main_multiply1785  instR291 (zll_main_multiply1785_inR72[128:1], zll_main_multiply1785_inR72[0], zll_main_multiply1785_outR72);
  assign zll_main_multiply603_in = {zll_main_multiply268_in[127:0], zll_main_multiply268_in[255:128], zll_main_multiply1785_outR72};
  assign id_inR219 = zll_main_multiply603_in[255:128];
  assign zll_main_multiply55_in = {zll_main_multiply603_in[127:0], zll_main_multiply603_in[383:256], zll_main_multiply603_in[255:128], id_inR219[54]};
  assign id_inR220 = zll_main_multiply55_in[128:1];
  assign zll_main_multiply1792_inR73 = {zll_main_multiply55_in[256:129], id_inR220[54]};
  ZLL_Main_multiply1792  instR292 (zll_main_multiply1792_inR73[128:1], zll_main_multiply1792_inR73[0], zll_main_multiply1792_outR73);
  assign zll_main_multiply1788_inR38 = {zll_main_multiply55_in[384:257], zll_main_multiply55_in[256:129], zll_main_multiply55_in[0]};
  ZLL_Main_multiply1788  instR293 (zll_main_multiply1788_inR38[256:129], zll_main_multiply1788_inR38[128:1], zll_main_multiply1788_outR38);
  assign zll_main_multiply23_in = {zll_main_multiply603_in[127:0], zll_main_multiply603_in[255:128], (zll_main_multiply1788_inR38[0] == 1'h1) ? zll_main_multiply1788_outR38 : zll_main_multiply1792_outR73};
  assign id_inR221 = zll_main_multiply23_in[383:256];
  assign rewire_prelude_not_inR73 = id_inR221[0];
  ReWire_Prelude_not  instR294 (rewire_prelude_not_inR73[0], rewire_prelude_not_outR73);
  assign zll_main_multiply1785_inR73 = {zll_main_multiply23_in[383:256], rewire_prelude_not_outR73};
  ZLL_Main_multiply1785  instR295 (zll_main_multiply1785_inR73[128:1], zll_main_multiply1785_inR73[0], zll_main_multiply1785_outR73);
  assign zll_main_multiply1399_in = {zll_main_multiply23_in[127:0], zll_main_multiply23_in[255:128], zll_main_multiply1785_outR73};
  assign id_inR222 = zll_main_multiply1399_in[255:128];
  assign zll_main_multiply1637_in = {zll_main_multiply1399_in[127:0], zll_main_multiply1399_in[383:256], zll_main_multiply1399_in[255:128], id_inR222[53]};
  assign id_inR223 = zll_main_multiply1637_in[128:1];
  assign zll_main_multiply1792_inR74 = {zll_main_multiply1637_in[256:129], id_inR223[53]};
  ZLL_Main_multiply1792  instR296 (zll_main_multiply1792_inR74[128:1], zll_main_multiply1792_inR74[0], zll_main_multiply1792_outR74);
  assign zll_main_multiply1788_inR39 = {zll_main_multiply1637_in[384:257], zll_main_multiply1637_in[256:129], zll_main_multiply1637_in[0]};
  ZLL_Main_multiply1788  instR297 (zll_main_multiply1788_inR39[256:129], zll_main_multiply1788_inR39[128:1], zll_main_multiply1788_outR39);
  assign zll_main_multiply1662_in = {zll_main_multiply1399_in[127:0], zll_main_multiply1399_in[255:128], (zll_main_multiply1788_inR39[0] == 1'h1) ? zll_main_multiply1788_outR39 : zll_main_multiply1792_outR74};
  assign id_inR224 = zll_main_multiply1662_in[383:256];
  assign rewire_prelude_not_inR74 = id_inR224[0];
  ReWire_Prelude_not  instR298 (rewire_prelude_not_inR74[0], rewire_prelude_not_outR74);
  assign zll_main_multiply1785_inR74 = {zll_main_multiply1662_in[383:256], rewire_prelude_not_outR74};
  ZLL_Main_multiply1785  instR299 (zll_main_multiply1785_inR74[128:1], zll_main_multiply1785_inR74[0], zll_main_multiply1785_outR74);
  assign zll_main_multiply1106_in = {zll_main_multiply1662_in[255:128], zll_main_multiply1662_in[127:0], zll_main_multiply1785_outR74};
  assign id_inR225 = zll_main_multiply1106_in[383:256];
  assign zll_main_multiply1264_in = {zll_main_multiply1106_in[383:256], zll_main_multiply1106_in[127:0], zll_main_multiply1106_in[255:128], id_inR225[52]};
  assign id_inR226 = zll_main_multiply1264_in[384:257];
  assign zll_main_multiply1792_inR75 = {zll_main_multiply1264_in[128:1], id_inR226[52]};
  ZLL_Main_multiply1792  instR300 (zll_main_multiply1792_inR75[128:1], zll_main_multiply1792_inR75[0], zll_main_multiply1792_outR75);
  assign zll_main_multiply1788_inR40 = {zll_main_multiply1264_in[256:129], zll_main_multiply1264_in[128:1], zll_main_multiply1264_in[0]};
  ZLL_Main_multiply1788  instR301 (zll_main_multiply1788_inR40[256:129], zll_main_multiply1788_inR40[128:1], zll_main_multiply1788_outR40);
  assign zll_main_multiply24_in = {zll_main_multiply1106_in[383:256], zll_main_multiply1106_in[127:0], (zll_main_multiply1788_inR40[0] == 1'h1) ? zll_main_multiply1788_outR40 : zll_main_multiply1792_outR75};
  assign id_inR227 = zll_main_multiply24_in[255:128];
  assign rewire_prelude_not_inR75 = id_inR227[0];
  ReWire_Prelude_not  instR302 (rewire_prelude_not_inR75[0], rewire_prelude_not_outR75);
  assign zll_main_multiply1785_inR75 = {zll_main_multiply24_in[255:128], rewire_prelude_not_outR75};
  ZLL_Main_multiply1785  instR303 (zll_main_multiply1785_inR75[128:1], zll_main_multiply1785_inR75[0], zll_main_multiply1785_outR75);
  assign zll_main_multiply172_in = {zll_main_multiply24_in[383:256], zll_main_multiply24_in[127:0], zll_main_multiply1785_outR75};
  assign id_inR228 = zll_main_multiply172_in[383:256];
  assign zll_main_multiply771_in = {zll_main_multiply172_in[127:0], zll_main_multiply172_in[383:256], zll_main_multiply172_in[255:128], id_inR228[51]};
  assign id_inR229 = zll_main_multiply771_in[256:129];
  assign zll_main_multiply1792_inR76 = {zll_main_multiply771_in[128:1], id_inR229[51]};
  ZLL_Main_multiply1792  instR304 (zll_main_multiply1792_inR76[128:1], zll_main_multiply1792_inR76[0], zll_main_multiply1792_outR76);
  assign zll_main_multiply1788_inR41 = {zll_main_multiply771_in[384:257], zll_main_multiply771_in[128:1], zll_main_multiply771_in[0]};
  ZLL_Main_multiply1788  instR305 (zll_main_multiply1788_inR41[256:129], zll_main_multiply1788_inR41[128:1], zll_main_multiply1788_outR41);
  assign zll_main_multiply1587_in = {zll_main_multiply172_in[127:0], zll_main_multiply172_in[383:256], (zll_main_multiply1788_inR41[0] == 1'h1) ? zll_main_multiply1788_outR41 : zll_main_multiply1792_outR76};
  assign id_inR230 = zll_main_multiply1587_in[383:256];
  assign rewire_prelude_not_inR76 = id_inR230[0];
  ReWire_Prelude_not  instR306 (rewire_prelude_not_inR76[0], rewire_prelude_not_outR76);
  assign zll_main_multiply1785_inR76 = {zll_main_multiply1587_in[383:256], rewire_prelude_not_outR76};
  ZLL_Main_multiply1785  instR307 (zll_main_multiply1785_inR76[128:1], zll_main_multiply1785_inR76[0], zll_main_multiply1785_outR76);
  assign zll_main_multiply1550_in = {zll_main_multiply1587_in[255:128], zll_main_multiply1587_in[127:0], zll_main_multiply1785_outR76};
  assign id_inR231 = zll_main_multiply1550_in[383:256];
  assign zll_main_multiply1167_in = {zll_main_multiply1550_in[127:0], zll_main_multiply1550_in[383:256], zll_main_multiply1550_in[255:128], id_inR231[50]};
  assign id_inR232 = zll_main_multiply1167_in[256:129];
  assign zll_main_multiply1792_inR77 = {zll_main_multiply1167_in[128:1], id_inR232[50]};
  ZLL_Main_multiply1792  instR308 (zll_main_multiply1792_inR77[128:1], zll_main_multiply1792_inR77[0], zll_main_multiply1792_outR77);
  assign zll_main_multiply1788_inR42 = {zll_main_multiply1167_in[384:257], zll_main_multiply1167_in[128:1], zll_main_multiply1167_in[0]};
  ZLL_Main_multiply1788  instR309 (zll_main_multiply1788_inR42[256:129], zll_main_multiply1788_inR42[128:1], zll_main_multiply1788_outR42);
  assign zll_main_multiply1251_in = {zll_main_multiply1550_in[127:0], zll_main_multiply1550_in[383:256], (zll_main_multiply1788_inR42[0] == 1'h1) ? zll_main_multiply1788_outR42 : zll_main_multiply1792_outR77};
  assign id_inR233 = zll_main_multiply1251_in[383:256];
  assign rewire_prelude_not_inR77 = id_inR233[0];
  ReWire_Prelude_not  instR310 (rewire_prelude_not_inR77[0], rewire_prelude_not_outR77);
  assign zll_main_multiply1785_inR77 = {zll_main_multiply1251_in[383:256], rewire_prelude_not_outR77};
  ZLL_Main_multiply1785  instR311 (zll_main_multiply1785_inR77[128:1], zll_main_multiply1785_inR77[0], zll_main_multiply1785_outR77);
  assign zll_main_multiply1320_in = {zll_main_multiply1251_in[255:128], zll_main_multiply1251_in[127:0], zll_main_multiply1785_outR77};
  assign id_inR234 = zll_main_multiply1320_in[383:256];
  assign zll_main_multiply43_in = {zll_main_multiply1320_in[127:0], zll_main_multiply1320_in[383:256], zll_main_multiply1320_in[255:128], id_inR234[49]};
  assign id_inR235 = zll_main_multiply43_in[256:129];
  assign zll_main_multiply1792_inR78 = {zll_main_multiply43_in[128:1], id_inR235[49]};
  ZLL_Main_multiply1792  instR312 (zll_main_multiply1792_inR78[128:1], zll_main_multiply1792_inR78[0], zll_main_multiply1792_outR78);
  assign zll_main_multiply1788_inR43 = {zll_main_multiply43_in[384:257], zll_main_multiply43_in[128:1], zll_main_multiply43_in[0]};
  ZLL_Main_multiply1788  instR313 (zll_main_multiply1788_inR43[256:129], zll_main_multiply1788_inR43[128:1], zll_main_multiply1788_outR43);
  assign zll_main_multiply1554_in = {zll_main_multiply1320_in[127:0], zll_main_multiply1320_in[383:256], (zll_main_multiply1788_inR43[0] == 1'h1) ? zll_main_multiply1788_outR43 : zll_main_multiply1792_outR78};
  assign id_inR236 = zll_main_multiply1554_in[383:256];
  assign rewire_prelude_not_inR78 = id_inR236[0];
  ReWire_Prelude_not  instR314 (rewire_prelude_not_inR78[0], rewire_prelude_not_outR78);
  assign zll_main_multiply1785_inR78 = {zll_main_multiply1554_in[383:256], rewire_prelude_not_outR78};
  ZLL_Main_multiply1785  instR315 (zll_main_multiply1785_inR78[128:1], zll_main_multiply1785_inR78[0], zll_main_multiply1785_outR78);
  assign zll_main_multiply257_in = {zll_main_multiply1554_in[127:0], zll_main_multiply1554_in[255:128], zll_main_multiply1785_outR78};
  assign id_inR237 = zll_main_multiply257_in[255:128];
  assign zll_main_multiply1513_in = {zll_main_multiply257_in[127:0], zll_main_multiply257_in[383:256], zll_main_multiply257_in[255:128], id_inR237[48]};
  assign id_inR238 = zll_main_multiply1513_in[128:1];
  assign zll_main_multiply1792_inR79 = {zll_main_multiply1513_in[256:129], id_inR238[48]};
  ZLL_Main_multiply1792  instR316 (zll_main_multiply1792_inR79[128:1], zll_main_multiply1792_inR79[0], zll_main_multiply1792_outR79);
  assign zll_main_multiply1788_inR44 = {zll_main_multiply1513_in[384:257], zll_main_multiply1513_in[256:129], zll_main_multiply1513_in[0]};
  ZLL_Main_multiply1788  instR317 (zll_main_multiply1788_inR44[256:129], zll_main_multiply1788_inR44[128:1], zll_main_multiply1788_outR44);
  assign zll_main_multiply113_in = {zll_main_multiply257_in[127:0], zll_main_multiply257_in[255:128], (zll_main_multiply1788_inR44[0] == 1'h1) ? zll_main_multiply1788_outR44 : zll_main_multiply1792_outR79};
  assign id_inR239 = zll_main_multiply113_in[383:256];
  assign rewire_prelude_not_inR79 = id_inR239[0];
  ReWire_Prelude_not  instR318 (rewire_prelude_not_inR79[0], rewire_prelude_not_outR79);
  assign zll_main_multiply1785_inR79 = {zll_main_multiply113_in[383:256], rewire_prelude_not_outR79};
  ZLL_Main_multiply1785  instR319 (zll_main_multiply1785_inR79[128:1], zll_main_multiply1785_inR79[0], zll_main_multiply1785_outR79);
  assign zll_main_multiply1091_in = {zll_main_multiply113_in[255:128], zll_main_multiply113_in[127:0], zll_main_multiply1785_outR79};
  assign id_inR240 = zll_main_multiply1091_in[383:256];
  assign zll_main_multiply1266_in = {zll_main_multiply1091_in[383:256], zll_main_multiply1091_in[127:0], zll_main_multiply1091_in[255:128], id_inR240[47]};
  assign id_inR241 = zll_main_multiply1266_in[384:257];
  assign zll_main_multiply1792_inR80 = {zll_main_multiply1266_in[128:1], id_inR241[47]};
  ZLL_Main_multiply1792  instR320 (zll_main_multiply1792_inR80[128:1], zll_main_multiply1792_inR80[0], zll_main_multiply1792_outR80);
  assign zll_main_multiply1788_inR45 = {zll_main_multiply1266_in[256:129], zll_main_multiply1266_in[128:1], zll_main_multiply1266_in[0]};
  ZLL_Main_multiply1788  instR321 (zll_main_multiply1788_inR45[256:129], zll_main_multiply1788_inR45[128:1], zll_main_multiply1788_outR45);
  assign zll_main_multiply418_in = {zll_main_multiply1091_in[383:256], zll_main_multiply1091_in[127:0], (zll_main_multiply1788_inR45[0] == 1'h1) ? zll_main_multiply1788_outR45 : zll_main_multiply1792_outR80};
  assign id_inR242 = zll_main_multiply418_in[255:128];
  assign rewire_prelude_not_inR80 = id_inR242[0];
  ReWire_Prelude_not  instR322 (rewire_prelude_not_inR80[0], rewire_prelude_not_outR80);
  assign zll_main_multiply1785_inR80 = {zll_main_multiply418_in[255:128], rewire_prelude_not_outR80};
  ZLL_Main_multiply1785  instR323 (zll_main_multiply1785_inR80[128:1], zll_main_multiply1785_inR80[0], zll_main_multiply1785_outR80);
  assign zll_main_multiply409_in = {zll_main_multiply418_in[383:256], zll_main_multiply418_in[127:0], zll_main_multiply1785_outR80};
  assign id_inR243 = zll_main_multiply409_in[383:256];
  assign zll_main_multiply726_in = {zll_main_multiply409_in[127:0], zll_main_multiply409_in[383:256], zll_main_multiply409_in[255:128], id_inR243[46]};
  assign id_inR244 = zll_main_multiply726_in[256:129];
  assign zll_main_multiply1792_inR81 = {zll_main_multiply726_in[128:1], id_inR244[46]};
  ZLL_Main_multiply1792  instR324 (zll_main_multiply1792_inR81[128:1], zll_main_multiply1792_inR81[0], zll_main_multiply1792_outR81);
  assign zll_main_multiply1788_inR46 = {zll_main_multiply726_in[384:257], zll_main_multiply726_in[128:1], zll_main_multiply726_in[0]};
  ZLL_Main_multiply1788  instR325 (zll_main_multiply1788_inR46[256:129], zll_main_multiply1788_inR46[128:1], zll_main_multiply1788_outR46);
  assign zll_main_multiply1387_in = {zll_main_multiply409_in[127:0], zll_main_multiply409_in[383:256], (zll_main_multiply1788_inR46[0] == 1'h1) ? zll_main_multiply1788_outR46 : zll_main_multiply1792_outR81};
  assign id_inR245 = zll_main_multiply1387_in[383:256];
  assign rewire_prelude_not_inR81 = id_inR245[0];
  ReWire_Prelude_not  instR326 (rewire_prelude_not_inR81[0], rewire_prelude_not_outR81);
  assign zll_main_multiply1785_inR81 = {zll_main_multiply1387_in[383:256], rewire_prelude_not_outR81};
  ZLL_Main_multiply1785  instR327 (zll_main_multiply1785_inR81[128:1], zll_main_multiply1785_inR81[0], zll_main_multiply1785_outR81);
  assign zll_main_multiply584_in = {zll_main_multiply1387_in[127:0], zll_main_multiply1387_in[255:128], zll_main_multiply1785_outR81};
  assign id_inR246 = zll_main_multiply584_in[255:128];
  assign zll_main_multiply764_in = {zll_main_multiply584_in[127:0], zll_main_multiply584_in[383:256], zll_main_multiply584_in[255:128], id_inR246[45]};
  assign id_inR247 = zll_main_multiply764_in[128:1];
  assign zll_main_multiply1792_inR82 = {zll_main_multiply764_in[256:129], id_inR247[45]};
  ZLL_Main_multiply1792  instR328 (zll_main_multiply1792_inR82[128:1], zll_main_multiply1792_inR82[0], zll_main_multiply1792_outR82);
  assign zll_main_multiply1788_inR47 = {zll_main_multiply764_in[384:257], zll_main_multiply764_in[256:129], zll_main_multiply764_in[0]};
  ZLL_Main_multiply1788  instR329 (zll_main_multiply1788_inR47[256:129], zll_main_multiply1788_inR47[128:1], zll_main_multiply1788_outR47);
  assign zll_main_multiply1627_in = {zll_main_multiply584_in[127:0], zll_main_multiply584_in[255:128], (zll_main_multiply1788_inR47[0] == 1'h1) ? zll_main_multiply1788_outR47 : zll_main_multiply1792_outR82};
  assign id_inR248 = zll_main_multiply1627_in[383:256];
  assign rewire_prelude_not_inR82 = id_inR248[0];
  ReWire_Prelude_not  instR330 (rewire_prelude_not_inR82[0], rewire_prelude_not_outR82);
  assign zll_main_multiply1785_inR82 = {zll_main_multiply1627_in[383:256], rewire_prelude_not_outR82};
  ZLL_Main_multiply1785  instR331 (zll_main_multiply1785_inR82[128:1], zll_main_multiply1785_inR82[0], zll_main_multiply1785_outR82);
  assign zll_main_multiply442_in = {zll_main_multiply1627_in[255:128], zll_main_multiply1627_in[127:0], zll_main_multiply1785_outR82};
  assign id_inR249 = zll_main_multiply442_in[383:256];
  assign zll_main_multiply1121_in = {zll_main_multiply442_in[127:0], zll_main_multiply442_in[383:256], zll_main_multiply442_in[255:128], id_inR249[44]};
  assign id_inR250 = zll_main_multiply1121_in[256:129];
  assign zll_main_multiply1792_inR83 = {zll_main_multiply1121_in[128:1], id_inR250[44]};
  ZLL_Main_multiply1792  instR332 (zll_main_multiply1792_inR83[128:1], zll_main_multiply1792_inR83[0], zll_main_multiply1792_outR83);
  assign zll_main_multiply1788_inR48 = {zll_main_multiply1121_in[384:257], zll_main_multiply1121_in[128:1], zll_main_multiply1121_in[0]};
  ZLL_Main_multiply1788  instR333 (zll_main_multiply1788_inR48[256:129], zll_main_multiply1788_inR48[128:1], zll_main_multiply1788_outR48);
  assign zll_main_multiply223_in = {zll_main_multiply442_in[127:0], zll_main_multiply442_in[383:256], (zll_main_multiply1788_inR48[0] == 1'h1) ? zll_main_multiply1788_outR48 : zll_main_multiply1792_outR83};
  assign id_inR251 = zll_main_multiply223_in[383:256];
  assign rewire_prelude_not_inR83 = id_inR251[0];
  ReWire_Prelude_not  instR334 (rewire_prelude_not_inR83[0], rewire_prelude_not_outR83);
  assign zll_main_multiply1785_inR83 = {zll_main_multiply223_in[383:256], rewire_prelude_not_outR83};
  ZLL_Main_multiply1785  instR335 (zll_main_multiply1785_inR83[128:1], zll_main_multiply1785_inR83[0], zll_main_multiply1785_outR83);
  assign zll_main_multiply1410_in = {zll_main_multiply223_in[255:128], zll_main_multiply223_in[127:0], zll_main_multiply1785_outR83};
  assign id_inR252 = zll_main_multiply1410_in[383:256];
  assign zll_main_multiply1147_in = {zll_main_multiply1410_in[127:0], zll_main_multiply1410_in[383:256], zll_main_multiply1410_in[255:128], id_inR252[43]};
  assign id_inR253 = zll_main_multiply1147_in[256:129];
  assign zll_main_multiply1792_inR84 = {zll_main_multiply1147_in[128:1], id_inR253[43]};
  ZLL_Main_multiply1792  instR336 (zll_main_multiply1792_inR84[128:1], zll_main_multiply1792_inR84[0], zll_main_multiply1792_outR84);
  assign zll_main_multiply1788_inR49 = {zll_main_multiply1147_in[384:257], zll_main_multiply1147_in[128:1], zll_main_multiply1147_in[0]};
  ZLL_Main_multiply1788  instR337 (zll_main_multiply1788_inR49[256:129], zll_main_multiply1788_inR49[128:1], zll_main_multiply1788_outR49);
  assign zll_main_multiply1137_in = {zll_main_multiply1410_in[127:0], zll_main_multiply1410_in[383:256], (zll_main_multiply1788_inR49[0] == 1'h1) ? zll_main_multiply1788_outR49 : zll_main_multiply1792_outR84};
  assign id_inR254 = zll_main_multiply1137_in[383:256];
  assign rewire_prelude_not_inR84 = id_inR254[0];
  ReWire_Prelude_not  instR338 (rewire_prelude_not_inR84[0], rewire_prelude_not_outR84);
  assign zll_main_multiply1785_inR84 = {zll_main_multiply1137_in[383:256], rewire_prelude_not_outR84};
  ZLL_Main_multiply1785  instR339 (zll_main_multiply1785_inR84[128:1], zll_main_multiply1785_inR84[0], zll_main_multiply1785_outR84);
  assign zll_main_multiply1582_in = {zll_main_multiply1137_in[127:0], zll_main_multiply1137_in[255:128], zll_main_multiply1785_outR84};
  assign id_inR255 = zll_main_multiply1582_in[255:128];
  assign zll_main_multiply47_in = {zll_main_multiply1582_in[383:256], zll_main_multiply1582_in[255:128], zll_main_multiply1582_in[127:0], id_inR255[42]};
  assign id_inR256 = zll_main_multiply47_in[256:129];
  assign zll_main_multiply1792_inR85 = {zll_main_multiply47_in[384:257], id_inR256[42]};
  ZLL_Main_multiply1792  instR340 (zll_main_multiply1792_inR85[128:1], zll_main_multiply1792_inR85[0], zll_main_multiply1792_outR85);
  assign zll_main_multiply1749_inR35 = {zll_main_multiply47_in[384:257], zll_main_multiply47_in[128:1], zll_main_multiply47_in[0]};
  ZLL_Main_multiply1749  instR341 (zll_main_multiply1749_inR35[256:129], zll_main_multiply1749_inR35[128:1], zll_main_multiply1749_outR35);
  assign zll_main_multiply1047_in = {zll_main_multiply1582_in[255:128], zll_main_multiply1582_in[127:0], (zll_main_multiply1749_inR35[0] == 1'h1) ? zll_main_multiply1749_outR35 : zll_main_multiply1792_outR85};
  assign id_inR257 = zll_main_multiply1047_in[255:128];
  assign rewire_prelude_not_inR85 = id_inR257[0];
  ReWire_Prelude_not  instR342 (rewire_prelude_not_inR85[0], rewire_prelude_not_outR85);
  assign zll_main_multiply1785_inR85 = {zll_main_multiply1047_in[255:128], rewire_prelude_not_outR85};
  ZLL_Main_multiply1785  instR343 (zll_main_multiply1785_inR85[128:1], zll_main_multiply1785_inR85[0], zll_main_multiply1785_outR85);
  assign zll_main_multiply98_in = {zll_main_multiply1047_in[127:0], zll_main_multiply1047_in[383:256], zll_main_multiply1785_outR85};
  assign id_inR258 = zll_main_multiply98_in[255:128];
  assign zll_main_multiply1104_in = {zll_main_multiply98_in[383:256], zll_main_multiply98_in[127:0], zll_main_multiply98_in[255:128], id_inR258[41]};
  assign id_inR259 = zll_main_multiply1104_in[128:1];
  assign zll_main_multiply1792_inR86 = {zll_main_multiply1104_in[384:257], id_inR259[41]};
  ZLL_Main_multiply1792  instR344 (zll_main_multiply1792_inR86[128:1], zll_main_multiply1792_inR86[0], zll_main_multiply1792_outR86);
  assign zll_main_multiply1749_inR36 = {zll_main_multiply1104_in[384:257], zll_main_multiply1104_in[256:129], zll_main_multiply1104_in[0]};
  ZLL_Main_multiply1749  instR345 (zll_main_multiply1749_inR36[256:129], zll_main_multiply1749_inR36[128:1], zll_main_multiply1749_outR36);
  assign zll_main_multiply345_in = {zll_main_multiply98_in[127:0], zll_main_multiply98_in[255:128], (zll_main_multiply1749_inR36[0] == 1'h1) ? zll_main_multiply1749_outR36 : zll_main_multiply1792_outR86};
  assign id_inR260 = zll_main_multiply345_in[383:256];
  assign rewire_prelude_not_inR86 = id_inR260[0];
  ReWire_Prelude_not  instR346 (rewire_prelude_not_inR86[0], rewire_prelude_not_outR86);
  assign zll_main_multiply1785_inR86 = {zll_main_multiply345_in[383:256], rewire_prelude_not_outR86};
  ZLL_Main_multiply1785  instR347 (zll_main_multiply1785_inR86[128:1], zll_main_multiply1785_inR86[0], zll_main_multiply1785_outR86);
  assign zll_main_multiply1438_in = {zll_main_multiply345_in[255:128], zll_main_multiply345_in[127:0], zll_main_multiply1785_outR86};
  assign id_inR261 = zll_main_multiply1438_in[383:256];
  assign zll_main_multiply1483_in = {zll_main_multiply1438_in[127:0], zll_main_multiply1438_in[383:256], zll_main_multiply1438_in[255:128], id_inR261[40]};
  assign id_inR262 = zll_main_multiply1483_in[256:129];
  assign zll_main_multiply1792_inR87 = {zll_main_multiply1483_in[128:1], id_inR262[40]};
  ZLL_Main_multiply1792  instR348 (zll_main_multiply1792_inR87[128:1], zll_main_multiply1792_inR87[0], zll_main_multiply1792_outR87);
  assign zll_main_multiply1788_inR50 = {zll_main_multiply1483_in[384:257], zll_main_multiply1483_in[128:1], zll_main_multiply1483_in[0]};
  ZLL_Main_multiply1788  instR349 (zll_main_multiply1788_inR50[256:129], zll_main_multiply1788_inR50[128:1], zll_main_multiply1788_outR50);
  assign zll_main_multiply56_in = {zll_main_multiply1438_in[127:0], zll_main_multiply1438_in[383:256], (zll_main_multiply1788_inR50[0] == 1'h1) ? zll_main_multiply1788_outR50 : zll_main_multiply1792_outR87};
  assign id_inR263 = zll_main_multiply56_in[383:256];
  assign rewire_prelude_not_inR87 = id_inR263[0];
  ReWire_Prelude_not  instR350 (rewire_prelude_not_inR87[0], rewire_prelude_not_outR87);
  assign zll_main_multiply1785_inR87 = {zll_main_multiply56_in[383:256], rewire_prelude_not_outR87};
  ZLL_Main_multiply1785  instR351 (zll_main_multiply1785_inR87[128:1], zll_main_multiply1785_inR87[0], zll_main_multiply1785_outR87);
  assign zll_main_multiply1200_in = {zll_main_multiply56_in[255:128], zll_main_multiply56_in[127:0], zll_main_multiply1785_outR87};
  assign id_inR264 = zll_main_multiply1200_in[383:256];
  assign zll_main_multiply800_in = {zll_main_multiply1200_in[127:0], zll_main_multiply1200_in[383:256], zll_main_multiply1200_in[255:128], id_inR264[39]};
  assign id_inR265 = zll_main_multiply800_in[256:129];
  assign zll_main_multiply1792_inR88 = {zll_main_multiply800_in[128:1], id_inR265[39]};
  ZLL_Main_multiply1792  instR352 (zll_main_multiply1792_inR88[128:1], zll_main_multiply1792_inR88[0], zll_main_multiply1792_outR88);
  assign zll_main_multiply1788_inR51 = {zll_main_multiply800_in[384:257], zll_main_multiply800_in[128:1], zll_main_multiply800_in[0]};
  ZLL_Main_multiply1788  instR353 (zll_main_multiply1788_inR51[256:129], zll_main_multiply1788_inR51[128:1], zll_main_multiply1788_outR51);
  assign zll_main_multiply411_in = {zll_main_multiply1200_in[127:0], zll_main_multiply1200_in[383:256], (zll_main_multiply1788_inR51[0] == 1'h1) ? zll_main_multiply1788_outR51 : zll_main_multiply1792_outR88};
  assign id_inR266 = zll_main_multiply411_in[383:256];
  assign rewire_prelude_not_inR88 = id_inR266[0];
  ReWire_Prelude_not  instR354 (rewire_prelude_not_inR88[0], rewire_prelude_not_outR88);
  assign zll_main_multiply1785_inR88 = {zll_main_multiply411_in[383:256], rewire_prelude_not_outR88};
  ZLL_Main_multiply1785  instR355 (zll_main_multiply1785_inR88[128:1], zll_main_multiply1785_inR88[0], zll_main_multiply1785_outR88);
  assign zll_main_multiply774_in = {zll_main_multiply411_in[255:128], zll_main_multiply411_in[127:0], zll_main_multiply1785_outR88};
  assign id_inR267 = zll_main_multiply774_in[383:256];
  assign zll_main_multiply129_in = {zll_main_multiply774_in[383:256], zll_main_multiply774_in[127:0], zll_main_multiply774_in[255:128], id_inR267[38]};
  assign id_inR268 = zll_main_multiply129_in[384:257];
  assign zll_main_multiply1792_inR89 = {zll_main_multiply129_in[128:1], id_inR268[38]};
  ZLL_Main_multiply1792  instR356 (zll_main_multiply1792_inR89[128:1], zll_main_multiply1792_inR89[0], zll_main_multiply1792_outR89);
  assign zll_main_multiply1788_inR52 = {zll_main_multiply129_in[256:129], zll_main_multiply129_in[128:1], zll_main_multiply129_in[0]};
  ZLL_Main_multiply1788  instR357 (zll_main_multiply1788_inR52[256:129], zll_main_multiply1788_inR52[128:1], zll_main_multiply1788_outR52);
  assign zll_main_multiply1583_in = {zll_main_multiply774_in[383:256], zll_main_multiply774_in[127:0], (zll_main_multiply1788_inR52[0] == 1'h1) ? zll_main_multiply1788_outR52 : zll_main_multiply1792_outR89};
  assign id_inR269 = zll_main_multiply1583_in[255:128];
  assign rewire_prelude_not_inR89 = id_inR269[0];
  ReWire_Prelude_not  instR358 (rewire_prelude_not_inR89[0], rewire_prelude_not_outR89);
  assign zll_main_multiply1785_inR89 = {zll_main_multiply1583_in[255:128], rewire_prelude_not_outR89};
  ZLL_Main_multiply1785  instR359 (zll_main_multiply1785_inR89[128:1], zll_main_multiply1785_inR89[0], zll_main_multiply1785_outR89);
  assign zll_main_multiply226_in = {zll_main_multiply1583_in[383:256], zll_main_multiply1583_in[127:0], zll_main_multiply1785_outR89};
  assign id_inR270 = zll_main_multiply226_in[383:256];
  assign zll_main_multiply434_in = {zll_main_multiply226_in[127:0], zll_main_multiply226_in[383:256], zll_main_multiply226_in[255:128], id_inR270[37]};
  assign id_inR271 = zll_main_multiply434_in[256:129];
  assign zll_main_multiply1792_inR90 = {zll_main_multiply434_in[128:1], id_inR271[37]};
  ZLL_Main_multiply1792  instR360 (zll_main_multiply1792_inR90[128:1], zll_main_multiply1792_inR90[0], zll_main_multiply1792_outR90);
  assign zll_main_multiply1788_inR53 = {zll_main_multiply434_in[384:257], zll_main_multiply434_in[128:1], zll_main_multiply434_in[0]};
  ZLL_Main_multiply1788  instR361 (zll_main_multiply1788_inR53[256:129], zll_main_multiply1788_inR53[128:1], zll_main_multiply1788_outR53);
  assign zll_main_multiply1369_in = {zll_main_multiply226_in[127:0], zll_main_multiply226_in[383:256], (zll_main_multiply1788_inR53[0] == 1'h1) ? zll_main_multiply1788_outR53 : zll_main_multiply1792_outR90};
  assign id_inR272 = zll_main_multiply1369_in[383:256];
  assign rewire_prelude_not_inR90 = id_inR272[0];
  ReWire_Prelude_not  instR362 (rewire_prelude_not_inR90[0], rewire_prelude_not_outR90);
  assign zll_main_multiply1785_inR90 = {zll_main_multiply1369_in[383:256], rewire_prelude_not_outR90};
  ZLL_Main_multiply1785  instR363 (zll_main_multiply1785_inR90[128:1], zll_main_multiply1785_inR90[0], zll_main_multiply1785_outR90);
  assign zll_main_multiply697_in = {zll_main_multiply1369_in[127:0], zll_main_multiply1369_in[255:128], zll_main_multiply1785_outR90};
  assign id_inR273 = zll_main_multiply697_in[255:128];
  assign zll_main_multiply869_in = {zll_main_multiply697_in[127:0], zll_main_multiply697_in[383:256], zll_main_multiply697_in[255:128], id_inR273[36]};
  assign id_inR274 = zll_main_multiply869_in[128:1];
  assign zll_main_multiply1792_inR91 = {zll_main_multiply869_in[256:129], id_inR274[36]};
  ZLL_Main_multiply1792  instR364 (zll_main_multiply1792_inR91[128:1], zll_main_multiply1792_inR91[0], zll_main_multiply1792_outR91);
  assign zll_main_multiply1788_inR54 = {zll_main_multiply869_in[384:257], zll_main_multiply869_in[256:129], zll_main_multiply869_in[0]};
  ZLL_Main_multiply1788  instR365 (zll_main_multiply1788_inR54[256:129], zll_main_multiply1788_inR54[128:1], zll_main_multiply1788_outR54);
  assign zll_main_multiply1774_in = {zll_main_multiply697_in[127:0], zll_main_multiply697_in[255:128], (zll_main_multiply1788_inR54[0] == 1'h1) ? zll_main_multiply1788_outR54 : zll_main_multiply1792_outR91};
  assign id_inR275 = zll_main_multiply1774_in[383:256];
  assign rewire_prelude_not_inR91 = id_inR275[0];
  ReWire_Prelude_not  instR366 (rewire_prelude_not_inR91[0], rewire_prelude_not_outR91);
  assign zll_main_multiply1785_inR91 = {zll_main_multiply1774_in[383:256], rewire_prelude_not_outR91};
  ZLL_Main_multiply1785  instR367 (zll_main_multiply1785_inR91[128:1], zll_main_multiply1785_inR91[0], zll_main_multiply1785_outR91);
  assign zll_main_multiply779_in = {zll_main_multiply1774_in[127:0], zll_main_multiply1774_in[255:128], zll_main_multiply1785_outR91};
  assign id_inR276 = zll_main_multiply779_in[255:128];
  assign zll_main_multiply1551_in = {zll_main_multiply779_in[383:256], zll_main_multiply779_in[255:128], zll_main_multiply779_in[127:0], id_inR276[35]};
  assign id_inR277 = zll_main_multiply1551_in[256:129];
  assign zll_main_multiply1792_inR92 = {zll_main_multiply1551_in[384:257], id_inR277[35]};
  ZLL_Main_multiply1792  instR368 (zll_main_multiply1792_inR92[128:1], zll_main_multiply1792_inR92[0], zll_main_multiply1792_outR92);
  assign zll_main_multiply1749_inR37 = {zll_main_multiply1551_in[384:257], zll_main_multiply1551_in[128:1], zll_main_multiply1551_in[0]};
  ZLL_Main_multiply1749  instR369 (zll_main_multiply1749_inR37[256:129], zll_main_multiply1749_inR37[128:1], zll_main_multiply1749_outR37);
  assign zll_main_multiply845_in = {zll_main_multiply779_in[255:128], zll_main_multiply779_in[127:0], (zll_main_multiply1749_inR37[0] == 1'h1) ? zll_main_multiply1749_outR37 : zll_main_multiply1792_outR92};
  assign id_inR278 = zll_main_multiply845_in[255:128];
  assign rewire_prelude_not_inR92 = id_inR278[0];
  ReWire_Prelude_not  instR370 (rewire_prelude_not_inR92[0], rewire_prelude_not_outR92);
  assign zll_main_multiply1785_inR92 = {zll_main_multiply845_in[255:128], rewire_prelude_not_outR92};
  ZLL_Main_multiply1785  instR371 (zll_main_multiply1785_inR92[128:1], zll_main_multiply1785_inR92[0], zll_main_multiply1785_outR92);
  assign zll_main_multiply565_in = {zll_main_multiply845_in[127:0], zll_main_multiply845_in[383:256], zll_main_multiply1785_outR92};
  assign id_inR279 = zll_main_multiply565_in[255:128];
  assign zll_main_multiply496_in = {zll_main_multiply565_in[127:0], zll_main_multiply565_in[383:256], zll_main_multiply565_in[255:128], id_inR279[34]};
  assign id_inR280 = zll_main_multiply496_in[128:1];
  assign zll_main_multiply1792_inR93 = {zll_main_multiply496_in[256:129], id_inR280[34]};
  ZLL_Main_multiply1792  instR372 (zll_main_multiply1792_inR93[128:1], zll_main_multiply1792_inR93[0], zll_main_multiply1792_outR93);
  assign zll_main_multiply1788_inR55 = {zll_main_multiply496_in[384:257], zll_main_multiply496_in[256:129], zll_main_multiply496_in[0]};
  ZLL_Main_multiply1788  instR373 (zll_main_multiply1788_inR55[256:129], zll_main_multiply1788_inR55[128:1], zll_main_multiply1788_outR55);
  assign zll_main_multiply1479_in = {zll_main_multiply565_in[127:0], zll_main_multiply565_in[255:128], (zll_main_multiply1788_inR55[0] == 1'h1) ? zll_main_multiply1788_outR55 : zll_main_multiply1792_outR93};
  assign id_inR281 = zll_main_multiply1479_in[383:256];
  assign rewire_prelude_not_inR93 = id_inR281[0];
  ReWire_Prelude_not  instR374 (rewire_prelude_not_inR93[0], rewire_prelude_not_outR93);
  assign zll_main_multiply1785_inR93 = {zll_main_multiply1479_in[383:256], rewire_prelude_not_outR93};
  ZLL_Main_multiply1785  instR375 (zll_main_multiply1785_inR93[128:1], zll_main_multiply1785_inR93[0], zll_main_multiply1785_outR93);
  assign zll_main_multiply703_in = {zll_main_multiply1479_in[127:0], zll_main_multiply1479_in[255:128], zll_main_multiply1785_outR93};
  assign id_inR282 = zll_main_multiply703_in[255:128];
  assign zll_main_multiply1286_in = {zll_main_multiply703_in[383:256], zll_main_multiply703_in[127:0], zll_main_multiply703_in[255:128], id_inR282[33]};
  assign id_inR283 = zll_main_multiply1286_in[128:1];
  assign zll_main_multiply1792_inR94 = {zll_main_multiply1286_in[384:257], id_inR283[33]};
  ZLL_Main_multiply1792  instR376 (zll_main_multiply1792_inR94[128:1], zll_main_multiply1792_inR94[0], zll_main_multiply1792_outR94);
  assign zll_main_multiply1749_inR38 = {zll_main_multiply1286_in[384:257], zll_main_multiply1286_in[256:129], zll_main_multiply1286_in[0]};
  ZLL_Main_multiply1749  instR377 (zll_main_multiply1749_inR38[256:129], zll_main_multiply1749_inR38[128:1], zll_main_multiply1749_outR38);
  assign zll_main_multiply293_in = {zll_main_multiply703_in[127:0], zll_main_multiply703_in[255:128], (zll_main_multiply1749_inR38[0] == 1'h1) ? zll_main_multiply1749_outR38 : zll_main_multiply1792_outR94};
  assign id_inR284 = zll_main_multiply293_in[383:256];
  assign rewire_prelude_not_inR94 = id_inR284[0];
  ReWire_Prelude_not  instR378 (rewire_prelude_not_inR94[0], rewire_prelude_not_outR94);
  assign zll_main_multiply1785_inR94 = {zll_main_multiply293_in[383:256], rewire_prelude_not_outR94};
  ZLL_Main_multiply1785  instR379 (zll_main_multiply1785_inR94[128:1], zll_main_multiply1785_inR94[0], zll_main_multiply1785_outR94);
  assign zll_main_multiply1290_in = {zll_main_multiply293_in[127:0], zll_main_multiply293_in[255:128], zll_main_multiply1785_outR94};
  assign id_inR285 = zll_main_multiply1290_in[255:128];
  assign zll_main_multiply1189_in = {zll_main_multiply1290_in[127:0], zll_main_multiply1290_in[383:256], zll_main_multiply1290_in[255:128], id_inR285[32]};
  assign id_inR286 = zll_main_multiply1189_in[128:1];
  assign zll_main_multiply1792_inR95 = {zll_main_multiply1189_in[256:129], id_inR286[32]};
  ZLL_Main_multiply1792  instR380 (zll_main_multiply1792_inR95[128:1], zll_main_multiply1792_inR95[0], zll_main_multiply1792_outR95);
  assign zll_main_multiply1788_inR56 = {zll_main_multiply1189_in[384:257], zll_main_multiply1189_in[256:129], zll_main_multiply1189_in[0]};
  ZLL_Main_multiply1788  instR381 (zll_main_multiply1788_inR56[256:129], zll_main_multiply1788_inR56[128:1], zll_main_multiply1788_outR56);
  assign zll_main_multiply1404_in = {zll_main_multiply1290_in[127:0], zll_main_multiply1290_in[255:128], (zll_main_multiply1788_inR56[0] == 1'h1) ? zll_main_multiply1788_outR56 : zll_main_multiply1792_outR95};
  assign id_inR287 = zll_main_multiply1404_in[383:256];
  assign rewire_prelude_not_inR95 = id_inR287[0];
  ReWire_Prelude_not  instR382 (rewire_prelude_not_inR95[0], rewire_prelude_not_outR95);
  assign zll_main_multiply1785_inR95 = {zll_main_multiply1404_in[383:256], rewire_prelude_not_outR95};
  ZLL_Main_multiply1785  instR383 (zll_main_multiply1785_inR95[128:1], zll_main_multiply1785_inR95[0], zll_main_multiply1785_outR95);
  assign zll_main_multiply676_in = {zll_main_multiply1404_in[127:0], zll_main_multiply1404_in[255:128], zll_main_multiply1785_outR95};
  assign id_inR288 = zll_main_multiply676_in[255:128];
  assign zll_main_multiply1769_in = {zll_main_multiply676_in[127:0], zll_main_multiply676_in[383:256], zll_main_multiply676_in[255:128], id_inR288[31]};
  assign id_inR289 = zll_main_multiply1769_in[128:1];
  assign zll_main_multiply1792_inR96 = {zll_main_multiply1769_in[256:129], id_inR289[31]};
  ZLL_Main_multiply1792  instR384 (zll_main_multiply1792_inR96[128:1], zll_main_multiply1792_inR96[0], zll_main_multiply1792_outR96);
  assign zll_main_multiply1788_inR57 = {zll_main_multiply1769_in[384:257], zll_main_multiply1769_in[256:129], zll_main_multiply1769_in[0]};
  ZLL_Main_multiply1788  instR385 (zll_main_multiply1788_inR57[256:129], zll_main_multiply1788_inR57[128:1], zll_main_multiply1788_outR57);
  assign zll_main_multiply464_in = {zll_main_multiply676_in[127:0], zll_main_multiply676_in[255:128], (zll_main_multiply1788_inR57[0] == 1'h1) ? zll_main_multiply1788_outR57 : zll_main_multiply1792_outR96};
  assign id_inR290 = zll_main_multiply464_in[383:256];
  assign rewire_prelude_not_inR96 = id_inR290[0];
  ReWire_Prelude_not  instR386 (rewire_prelude_not_inR96[0], rewire_prelude_not_outR96);
  assign zll_main_multiply1785_inR96 = {zll_main_multiply464_in[383:256], rewire_prelude_not_outR96};
  ZLL_Main_multiply1785  instR387 (zll_main_multiply1785_inR96[128:1], zll_main_multiply1785_inR96[0], zll_main_multiply1785_outR96);
  assign zll_main_multiply538_in = {zll_main_multiply464_in[127:0], zll_main_multiply464_in[255:128], zll_main_multiply1785_outR96};
  assign id_inR291 = zll_main_multiply538_in[255:128];
  assign zll_main_multiply175_in = {zll_main_multiply538_in[383:256], zll_main_multiply538_in[127:0], zll_main_multiply538_in[255:128], id_inR291[30]};
  assign id_inR292 = zll_main_multiply175_in[128:1];
  assign zll_main_multiply1792_inR97 = {zll_main_multiply175_in[384:257], id_inR292[30]};
  ZLL_Main_multiply1792  instR388 (zll_main_multiply1792_inR97[128:1], zll_main_multiply1792_inR97[0], zll_main_multiply1792_outR97);
  assign zll_main_multiply1749_inR39 = {zll_main_multiply175_in[384:257], zll_main_multiply175_in[256:129], zll_main_multiply175_in[0]};
  ZLL_Main_multiply1749  instR389 (zll_main_multiply1749_inR39[256:129], zll_main_multiply1749_inR39[128:1], zll_main_multiply1749_outR39);
  assign zll_main_multiply376_in = {zll_main_multiply538_in[127:0], zll_main_multiply538_in[255:128], (zll_main_multiply1749_inR39[0] == 1'h1) ? zll_main_multiply1749_outR39 : zll_main_multiply1792_outR97};
  assign id_inR293 = zll_main_multiply376_in[383:256];
  assign rewire_prelude_not_inR97 = id_inR293[0];
  ReWire_Prelude_not  instR390 (rewire_prelude_not_inR97[0], rewire_prelude_not_outR97);
  assign zll_main_multiply1785_inR97 = {zll_main_multiply376_in[383:256], rewire_prelude_not_outR97};
  ZLL_Main_multiply1785  instR391 (zll_main_multiply1785_inR97[128:1], zll_main_multiply1785_inR97[0], zll_main_multiply1785_outR97);
  assign zll_main_multiply471_in = {zll_main_multiply376_in[127:0], zll_main_multiply376_in[255:128], zll_main_multiply1785_outR97};
  assign id_inR294 = zll_main_multiply471_in[255:128];
  assign zll_main_multiply872_in = {zll_main_multiply471_in[127:0], zll_main_multiply471_in[383:256], zll_main_multiply471_in[255:128], id_inR294[29]};
  assign id_inR295 = zll_main_multiply872_in[128:1];
  assign zll_main_multiply1792_inR98 = {zll_main_multiply872_in[256:129], id_inR295[29]};
  ZLL_Main_multiply1792  instR392 (zll_main_multiply1792_inR98[128:1], zll_main_multiply1792_inR98[0], zll_main_multiply1792_outR98);
  assign zll_main_multiply1788_inR58 = {zll_main_multiply872_in[384:257], zll_main_multiply872_in[256:129], zll_main_multiply872_in[0]};
  ZLL_Main_multiply1788  instR393 (zll_main_multiply1788_inR58[256:129], zll_main_multiply1788_inR58[128:1], zll_main_multiply1788_outR58);
  assign zll_main_multiply1031_in = {zll_main_multiply471_in[127:0], zll_main_multiply471_in[255:128], (zll_main_multiply1788_inR58[0] == 1'h1) ? zll_main_multiply1788_outR58 : zll_main_multiply1792_outR98};
  assign id_inR296 = zll_main_multiply1031_in[383:256];
  assign rewire_prelude_not_inR98 = id_inR296[0];
  ReWire_Prelude_not  instR394 (rewire_prelude_not_inR98[0], rewire_prelude_not_outR98);
  assign zll_main_multiply1785_inR98 = {zll_main_multiply1031_in[383:256], rewire_prelude_not_outR98};
  ZLL_Main_multiply1785  instR395 (zll_main_multiply1785_inR98[128:1], zll_main_multiply1785_inR98[0], zll_main_multiply1785_outR98);
  assign zll_main_multiply639_in = {zll_main_multiply1031_in[127:0], zll_main_multiply1031_in[255:128], zll_main_multiply1785_outR98};
  assign id_inR297 = zll_main_multiply639_in[255:128];
  assign zll_main_multiply401_in = {zll_main_multiply639_in[383:256], zll_main_multiply639_in[127:0], zll_main_multiply639_in[255:128], id_inR297[28]};
  assign id_inR298 = zll_main_multiply401_in[128:1];
  assign zll_main_multiply1792_inR99 = {zll_main_multiply401_in[384:257], id_inR298[28]};
  ZLL_Main_multiply1792  instR396 (zll_main_multiply1792_inR99[128:1], zll_main_multiply1792_inR99[0], zll_main_multiply1792_outR99);
  assign zll_main_multiply1749_inR40 = {zll_main_multiply401_in[384:257], zll_main_multiply401_in[256:129], zll_main_multiply401_in[0]};
  ZLL_Main_multiply1749  instR397 (zll_main_multiply1749_inR40[256:129], zll_main_multiply1749_inR40[128:1], zll_main_multiply1749_outR40);
  assign zll_main_multiply1588_in = {zll_main_multiply639_in[127:0], zll_main_multiply639_in[255:128], (zll_main_multiply1749_inR40[0] == 1'h1) ? zll_main_multiply1749_outR40 : zll_main_multiply1792_outR99};
  assign id_inR299 = zll_main_multiply1588_in[383:256];
  assign rewire_prelude_not_inR99 = id_inR299[0];
  ReWire_Prelude_not  instR398 (rewire_prelude_not_inR99[0], rewire_prelude_not_outR99);
  assign zll_main_multiply1785_inR99 = {zll_main_multiply1588_in[383:256], rewire_prelude_not_outR99};
  ZLL_Main_multiply1785  instR399 (zll_main_multiply1785_inR99[128:1], zll_main_multiply1785_inR99[0], zll_main_multiply1785_outR99);
  assign zll_main_multiply1029_in = {zll_main_multiply1588_in[127:0], zll_main_multiply1588_in[255:128], zll_main_multiply1785_outR99};
  assign id_inR300 = zll_main_multiply1029_in[255:128];
  assign zll_main_multiply1340_in = {zll_main_multiply1029_in[127:0], zll_main_multiply1029_in[383:256], zll_main_multiply1029_in[255:128], id_inR300[27]};
  assign id_inR301 = zll_main_multiply1340_in[128:1];
  assign zll_main_multiply1792_inR100 = {zll_main_multiply1340_in[256:129], id_inR301[27]};
  ZLL_Main_multiply1792  instR400 (zll_main_multiply1792_inR100[128:1], zll_main_multiply1792_inR100[0], zll_main_multiply1792_outR100);
  assign zll_main_multiply1788_inR59 = {zll_main_multiply1340_in[384:257], zll_main_multiply1340_in[256:129], zll_main_multiply1340_in[0]};
  ZLL_Main_multiply1788  instR401 (zll_main_multiply1788_inR59[256:129], zll_main_multiply1788_inR59[128:1], zll_main_multiply1788_outR59);
  assign zll_main_multiply1080_in = {zll_main_multiply1029_in[127:0], zll_main_multiply1029_in[255:128], (zll_main_multiply1788_inR59[0] == 1'h1) ? zll_main_multiply1788_outR59 : zll_main_multiply1792_outR100};
  assign id_inR302 = zll_main_multiply1080_in[383:256];
  assign rewire_prelude_not_inR100 = id_inR302[0];
  ReWire_Prelude_not  instR402 (rewire_prelude_not_inR100[0], rewire_prelude_not_outR100);
  assign zll_main_multiply1785_inR100 = {zll_main_multiply1080_in[383:256], rewire_prelude_not_outR100};
  ZLL_Main_multiply1785  instR403 (zll_main_multiply1785_inR100[128:1], zll_main_multiply1785_inR100[0], zll_main_multiply1785_outR100);
  assign zll_main_multiply988_in = {zll_main_multiply1080_in[127:0], zll_main_multiply1080_in[255:128], zll_main_multiply1785_outR100};
  assign id_inR303 = zll_main_multiply988_in[255:128];
  assign zll_main_multiply1510_in = {zll_main_multiply988_in[383:256], zll_main_multiply988_in[255:128], zll_main_multiply988_in[127:0], id_inR303[26]};
  assign id_inR304 = zll_main_multiply1510_in[256:129];
  assign zll_main_multiply1792_inR101 = {zll_main_multiply1510_in[384:257], id_inR304[26]};
  ZLL_Main_multiply1792  instR404 (zll_main_multiply1792_inR101[128:1], zll_main_multiply1792_inR101[0], zll_main_multiply1792_outR101);
  assign zll_main_multiply1749_inR41 = {zll_main_multiply1510_in[384:257], zll_main_multiply1510_in[128:1], zll_main_multiply1510_in[0]};
  ZLL_Main_multiply1749  instR405 (zll_main_multiply1749_inR41[256:129], zll_main_multiply1749_inR41[128:1], zll_main_multiply1749_outR41);
  assign zll_main_multiply137_in = {zll_main_multiply988_in[255:128], zll_main_multiply988_in[127:0], (zll_main_multiply1749_inR41[0] == 1'h1) ? zll_main_multiply1749_outR41 : zll_main_multiply1792_outR101};
  assign id_inR305 = zll_main_multiply137_in[255:128];
  assign rewire_prelude_not_inR101 = id_inR305[0];
  ReWire_Prelude_not  instR406 (rewire_prelude_not_inR101[0], rewire_prelude_not_outR101);
  assign zll_main_multiply1785_inR101 = {zll_main_multiply137_in[255:128], rewire_prelude_not_outR101};
  ZLL_Main_multiply1785  instR407 (zll_main_multiply1785_inR101[128:1], zll_main_multiply1785_inR101[0], zll_main_multiply1785_outR101);
  assign zll_main_multiply67_in = {zll_main_multiply137_in[127:0], zll_main_multiply137_in[383:256], zll_main_multiply1785_outR101};
  assign id_inR306 = zll_main_multiply67_in[255:128];
  assign zll_main_multiply1678_in = {zll_main_multiply67_in[127:0], zll_main_multiply67_in[383:256], zll_main_multiply67_in[255:128], id_inR306[25]};
  assign id_inR307 = zll_main_multiply1678_in[128:1];
  assign zll_main_multiply1792_inR102 = {zll_main_multiply1678_in[256:129], id_inR307[25]};
  ZLL_Main_multiply1792  instR408 (zll_main_multiply1792_inR102[128:1], zll_main_multiply1792_inR102[0], zll_main_multiply1792_outR102);
  assign zll_main_multiply1788_inR60 = {zll_main_multiply1678_in[384:257], zll_main_multiply1678_in[256:129], zll_main_multiply1678_in[0]};
  ZLL_Main_multiply1788  instR409 (zll_main_multiply1788_inR60[256:129], zll_main_multiply1788_inR60[128:1], zll_main_multiply1788_outR60);
  assign zll_main_multiply662_in = {zll_main_multiply67_in[127:0], zll_main_multiply67_in[255:128], (zll_main_multiply1788_inR60[0] == 1'h1) ? zll_main_multiply1788_outR60 : zll_main_multiply1792_outR102};
  assign id_inR308 = zll_main_multiply662_in[383:256];
  assign rewire_prelude_not_inR102 = id_inR308[0];
  ReWire_Prelude_not  instR410 (rewire_prelude_not_inR102[0], rewire_prelude_not_outR102);
  assign zll_main_multiply1785_inR102 = {zll_main_multiply662_in[383:256], rewire_prelude_not_outR102};
  ZLL_Main_multiply1785  instR411 (zll_main_multiply1785_inR102[128:1], zll_main_multiply1785_inR102[0], zll_main_multiply1785_outR102);
  assign zll_main_multiply319_in = {zll_main_multiply662_in[255:128], zll_main_multiply662_in[127:0], zll_main_multiply1785_outR102};
  assign id_inR309 = zll_main_multiply319_in[383:256];
  assign zll_main_multiply817_in = {zll_main_multiply319_in[383:256], zll_main_multiply319_in[255:128], zll_main_multiply319_in[127:0], id_inR309[24]};
  assign id_inR310 = zll_main_multiply817_in[384:257];
  assign zll_main_multiply1792_inR103 = {zll_main_multiply817_in[256:129], id_inR310[24]};
  ZLL_Main_multiply1792  instR412 (zll_main_multiply1792_inR103[128:1], zll_main_multiply1792_inR103[0], zll_main_multiply1792_outR103);
  assign zll_main_multiply1749_inR42 = {zll_main_multiply817_in[256:129], zll_main_multiply817_in[128:1], zll_main_multiply817_in[0]};
  ZLL_Main_multiply1749  instR413 (zll_main_multiply1749_inR42[256:129], zll_main_multiply1749_inR42[128:1], zll_main_multiply1749_outR42);
  assign zll_main_multiply2_in = {zll_main_multiply319_in[383:256], zll_main_multiply319_in[127:0], (zll_main_multiply1749_inR42[0] == 1'h1) ? zll_main_multiply1749_outR42 : zll_main_multiply1792_outR103};
  assign id_inR311 = zll_main_multiply2_in[255:128];
  assign rewire_prelude_not_inR103 = id_inR311[0];
  ReWire_Prelude_not  instR414 (rewire_prelude_not_inR103[0], rewire_prelude_not_outR103);
  assign zll_main_multiply1785_inR103 = {zll_main_multiply2_in[255:128], rewire_prelude_not_outR103};
  ZLL_Main_multiply1785  instR415 (zll_main_multiply1785_inR103[128:1], zll_main_multiply1785_inR103[0], zll_main_multiply1785_outR103);
  assign zll_main_multiply912_in = {zll_main_multiply2_in[127:0], zll_main_multiply2_in[383:256], zll_main_multiply1785_outR103};
  assign id_inR312 = zll_main_multiply912_in[255:128];
  assign zll_main_multiply1624_in = {zll_main_multiply912_in[383:256], zll_main_multiply912_in[255:128], zll_main_multiply912_in[127:0], id_inR312[23]};
  assign id_inR313 = zll_main_multiply1624_in[256:129];
  assign zll_main_multiply1792_inR104 = {zll_main_multiply1624_in[384:257], id_inR313[23]};
  ZLL_Main_multiply1792  instR416 (zll_main_multiply1792_inR104[128:1], zll_main_multiply1792_inR104[0], zll_main_multiply1792_outR104);
  assign zll_main_multiply1749_inR43 = {zll_main_multiply1624_in[384:257], zll_main_multiply1624_in[128:1], zll_main_multiply1624_in[0]};
  ZLL_Main_multiply1749  instR417 (zll_main_multiply1749_inR43[256:129], zll_main_multiply1749_inR43[128:1], zll_main_multiply1749_outR43);
  assign zll_main_multiply977_in = {zll_main_multiply912_in[255:128], zll_main_multiply912_in[127:0], (zll_main_multiply1749_inR43[0] == 1'h1) ? zll_main_multiply1749_outR43 : zll_main_multiply1792_outR104};
  assign id_inR314 = zll_main_multiply977_in[255:128];
  assign rewire_prelude_not_inR104 = id_inR314[0];
  ReWire_Prelude_not  instR418 (rewire_prelude_not_inR104[0], rewire_prelude_not_outR104);
  assign zll_main_multiply1785_inR104 = {zll_main_multiply977_in[255:128], rewire_prelude_not_outR104};
  ZLL_Main_multiply1785  instR419 (zll_main_multiply1785_inR104[128:1], zll_main_multiply1785_inR104[0], zll_main_multiply1785_outR104);
  assign zll_main_multiply180_in = {zll_main_multiply977_in[127:0], zll_main_multiply977_in[383:256], zll_main_multiply1785_outR104};
  assign id_inR315 = zll_main_multiply180_in[255:128];
  assign zll_main_multiply476_in = {zll_main_multiply180_in[383:256], zll_main_multiply180_in[255:128], zll_main_multiply180_in[127:0], id_inR315[22]};
  assign id_inR316 = zll_main_multiply476_in[256:129];
  assign zll_main_multiply1792_inR105 = {zll_main_multiply476_in[384:257], id_inR316[22]};
  ZLL_Main_multiply1792  instR420 (zll_main_multiply1792_inR105[128:1], zll_main_multiply1792_inR105[0], zll_main_multiply1792_outR105);
  assign zll_main_multiply1749_inR44 = {zll_main_multiply476_in[384:257], zll_main_multiply476_in[128:1], zll_main_multiply476_in[0]};
  ZLL_Main_multiply1749  instR421 (zll_main_multiply1749_inR44[256:129], zll_main_multiply1749_inR44[128:1], zll_main_multiply1749_outR44);
  assign zll_main_multiply1599_in = {zll_main_multiply180_in[255:128], zll_main_multiply180_in[127:0], (zll_main_multiply1749_inR44[0] == 1'h1) ? zll_main_multiply1749_outR44 : zll_main_multiply1792_outR105};
  assign id_inR317 = zll_main_multiply1599_in[255:128];
  assign rewire_prelude_not_inR105 = id_inR317[0];
  ReWire_Prelude_not  instR422 (rewire_prelude_not_inR105[0], rewire_prelude_not_outR105);
  assign zll_main_multiply1785_inR105 = {zll_main_multiply1599_in[255:128], rewire_prelude_not_outR105};
  ZLL_Main_multiply1785  instR423 (zll_main_multiply1785_inR105[128:1], zll_main_multiply1785_inR105[0], zll_main_multiply1785_outR105);
  assign zll_main_multiply255_in = {zll_main_multiply1599_in[127:0], zll_main_multiply1599_in[383:256], zll_main_multiply1785_outR105};
  assign id_inR318 = zll_main_multiply255_in[255:128];
  assign zll_main_multiply1531_in = {zll_main_multiply255_in[383:256], zll_main_multiply255_in[127:0], zll_main_multiply255_in[255:128], id_inR318[21]};
  assign id_inR319 = zll_main_multiply1531_in[128:1];
  assign zll_main_multiply1792_inR106 = {zll_main_multiply1531_in[384:257], id_inR319[21]};
  ZLL_Main_multiply1792  instR424 (zll_main_multiply1792_inR106[128:1], zll_main_multiply1792_inR106[0], zll_main_multiply1792_outR106);
  assign zll_main_multiply1749_inR45 = {zll_main_multiply1531_in[384:257], zll_main_multiply1531_in[256:129], zll_main_multiply1531_in[0]};
  ZLL_Main_multiply1749  instR425 (zll_main_multiply1749_inR45[256:129], zll_main_multiply1749_inR45[128:1], zll_main_multiply1749_outR45);
  assign zll_main_multiply1083_in = {zll_main_multiply255_in[127:0], zll_main_multiply255_in[255:128], (zll_main_multiply1749_inR45[0] == 1'h1) ? zll_main_multiply1749_outR45 : zll_main_multiply1792_outR106};
  assign id_inR320 = zll_main_multiply1083_in[383:256];
  assign rewire_prelude_not_inR106 = id_inR320[0];
  ReWire_Prelude_not  instR426 (rewire_prelude_not_inR106[0], rewire_prelude_not_outR106);
  assign zll_main_multiply1785_inR106 = {zll_main_multiply1083_in[383:256], rewire_prelude_not_outR106};
  ZLL_Main_multiply1785  instR427 (zll_main_multiply1785_inR106[128:1], zll_main_multiply1785_inR106[0], zll_main_multiply1785_outR106);
  assign zll_main_multiply989_in = {zll_main_multiply1083_in[127:0], zll_main_multiply1083_in[255:128], zll_main_multiply1785_outR106};
  assign id_inR321 = zll_main_multiply989_in[255:128];
  assign zll_main_multiply947_in = {zll_main_multiply989_in[383:256], zll_main_multiply989_in[127:0], zll_main_multiply989_in[255:128], id_inR321[20]};
  assign id_inR322 = zll_main_multiply947_in[128:1];
  assign zll_main_multiply1792_inR107 = {zll_main_multiply947_in[384:257], id_inR322[20]};
  ZLL_Main_multiply1792  instR428 (zll_main_multiply1792_inR107[128:1], zll_main_multiply1792_inR107[0], zll_main_multiply1792_outR107);
  assign zll_main_multiply1749_inR46 = {zll_main_multiply947_in[384:257], zll_main_multiply947_in[256:129], zll_main_multiply947_in[0]};
  ZLL_Main_multiply1749  instR429 (zll_main_multiply1749_inR46[256:129], zll_main_multiply1749_inR46[128:1], zll_main_multiply1749_outR46);
  assign zll_main_multiply1245_in = {zll_main_multiply989_in[127:0], zll_main_multiply989_in[255:128], (zll_main_multiply1749_inR46[0] == 1'h1) ? zll_main_multiply1749_outR46 : zll_main_multiply1792_outR107};
  assign id_inR323 = zll_main_multiply1245_in[383:256];
  assign rewire_prelude_not_inR107 = id_inR323[0];
  ReWire_Prelude_not  instR430 (rewire_prelude_not_inR107[0], rewire_prelude_not_outR107);
  assign zll_main_multiply1785_inR107 = {zll_main_multiply1245_in[383:256], rewire_prelude_not_outR107};
  ZLL_Main_multiply1785  instR431 (zll_main_multiply1785_inR107[128:1], zll_main_multiply1785_inR107[0], zll_main_multiply1785_outR107);
  assign zll_main_multiply167_in = {zll_main_multiply1245_in[127:0], zll_main_multiply1245_in[255:128], zll_main_multiply1785_outR107};
  assign id_inR324 = zll_main_multiply167_in[255:128];
  assign zll_main_multiply1045_in = {zll_main_multiply167_in[383:256], zll_main_multiply167_in[255:128], zll_main_multiply167_in[127:0], id_inR324[19]};
  assign id_inR325 = zll_main_multiply1045_in[256:129];
  assign zll_main_multiply1792_inR108 = {zll_main_multiply1045_in[384:257], id_inR325[19]};
  ZLL_Main_multiply1792  instR432 (zll_main_multiply1792_inR108[128:1], zll_main_multiply1792_inR108[0], zll_main_multiply1792_outR108);
  assign zll_main_multiply1749_inR47 = {zll_main_multiply1045_in[384:257], zll_main_multiply1045_in[128:1], zll_main_multiply1045_in[0]};
  ZLL_Main_multiply1749  instR433 (zll_main_multiply1749_inR47[256:129], zll_main_multiply1749_inR47[128:1], zll_main_multiply1749_outR47);
  assign zll_main_multiply348_in = {zll_main_multiply167_in[255:128], zll_main_multiply167_in[127:0], (zll_main_multiply1749_inR47[0] == 1'h1) ? zll_main_multiply1749_outR47 : zll_main_multiply1792_outR108};
  assign id_inR326 = zll_main_multiply348_in[255:128];
  assign rewire_prelude_not_inR108 = id_inR326[0];
  ReWire_Prelude_not  instR434 (rewire_prelude_not_inR108[0], rewire_prelude_not_outR108);
  assign zll_main_multiply1785_inR108 = {zll_main_multiply348_in[255:128], rewire_prelude_not_outR108};
  ZLL_Main_multiply1785  instR435 (zll_main_multiply1785_inR108[128:1], zll_main_multiply1785_inR108[0], zll_main_multiply1785_outR108);
  assign zll_main_multiply444_in = {zll_main_multiply348_in[127:0], zll_main_multiply348_in[383:256], zll_main_multiply1785_outR108};
  assign id_inR327 = zll_main_multiply444_in[255:128];
  assign zll_main_multiply19_in = {zll_main_multiply444_in[127:0], zll_main_multiply444_in[383:256], zll_main_multiply444_in[255:128], id_inR327[18]};
  assign id_inR328 = zll_main_multiply19_in[128:1];
  assign zll_main_multiply1792_inR109 = {zll_main_multiply19_in[256:129], id_inR328[18]};
  ZLL_Main_multiply1792  instR436 (zll_main_multiply1792_inR109[128:1], zll_main_multiply1792_inR109[0], zll_main_multiply1792_outR109);
  assign zll_main_multiply1788_inR61 = {zll_main_multiply19_in[384:257], zll_main_multiply19_in[256:129], zll_main_multiply19_in[0]};
  ZLL_Main_multiply1788  instR437 (zll_main_multiply1788_inR61[256:129], zll_main_multiply1788_inR61[128:1], zll_main_multiply1788_outR61);
  assign zll_main_multiply130_in = {zll_main_multiply444_in[127:0], zll_main_multiply444_in[255:128], (zll_main_multiply1788_inR61[0] == 1'h1) ? zll_main_multiply1788_outR61 : zll_main_multiply1792_outR109};
  assign id_inR329 = zll_main_multiply130_in[383:256];
  assign rewire_prelude_not_inR109 = id_inR329[0];
  ReWire_Prelude_not  instR438 (rewire_prelude_not_inR109[0], rewire_prelude_not_outR109);
  assign zll_main_multiply1785_inR109 = {zll_main_multiply130_in[383:256], rewire_prelude_not_outR109};
  ZLL_Main_multiply1785  instR439 (zll_main_multiply1785_inR109[128:1], zll_main_multiply1785_inR109[0], zll_main_multiply1785_outR109);
  assign zll_main_multiply1403_in = {zll_main_multiply130_in[127:0], zll_main_multiply130_in[255:128], zll_main_multiply1785_outR109};
  assign id_inR330 = zll_main_multiply1403_in[255:128];
  assign zll_main_multiply1323_in = {zll_main_multiply1403_in[383:256], zll_main_multiply1403_in[255:128], zll_main_multiply1403_in[127:0], id_inR330[17]};
  assign id_inR331 = zll_main_multiply1323_in[256:129];
  assign zll_main_multiply1792_inR110 = {zll_main_multiply1323_in[384:257], id_inR331[17]};
  ZLL_Main_multiply1792  instR440 (zll_main_multiply1792_inR110[128:1], zll_main_multiply1792_inR110[0], zll_main_multiply1792_outR110);
  assign zll_main_multiply1749_inR48 = {zll_main_multiply1323_in[384:257], zll_main_multiply1323_in[128:1], zll_main_multiply1323_in[0]};
  ZLL_Main_multiply1749  instR441 (zll_main_multiply1749_inR48[256:129], zll_main_multiply1749_inR48[128:1], zll_main_multiply1749_outR48);
  assign zll_main_multiply1329_in = {zll_main_multiply1403_in[255:128], zll_main_multiply1403_in[127:0], (zll_main_multiply1749_inR48[0] == 1'h1) ? zll_main_multiply1749_outR48 : zll_main_multiply1792_outR110};
  assign id_inR332 = zll_main_multiply1329_in[255:128];
  assign rewire_prelude_not_inR110 = id_inR332[0];
  ReWire_Prelude_not  instR442 (rewire_prelude_not_inR110[0], rewire_prelude_not_outR110);
  assign zll_main_multiply1785_inR110 = {zll_main_multiply1329_in[255:128], rewire_prelude_not_outR110};
  ZLL_Main_multiply1785  instR443 (zll_main_multiply1785_inR110[128:1], zll_main_multiply1785_inR110[0], zll_main_multiply1785_outR110);
  assign zll_main_multiply389_in = {zll_main_multiply1329_in[127:0], zll_main_multiply1329_in[383:256], zll_main_multiply1785_outR110};
  assign id_inR333 = zll_main_multiply389_in[255:128];
  assign zll_main_multiply294_in = {zll_main_multiply389_in[383:256], zll_main_multiply389_in[255:128], zll_main_multiply389_in[127:0], id_inR333[16]};
  assign id_inR334 = zll_main_multiply294_in[256:129];
  assign zll_main_multiply1792_inR111 = {zll_main_multiply294_in[384:257], id_inR334[16]};
  ZLL_Main_multiply1792  instR444 (zll_main_multiply1792_inR111[128:1], zll_main_multiply1792_inR111[0], zll_main_multiply1792_outR111);
  assign zll_main_multiply1749_inR49 = {zll_main_multiply294_in[384:257], zll_main_multiply294_in[128:1], zll_main_multiply294_in[0]};
  ZLL_Main_multiply1749  instR445 (zll_main_multiply1749_inR49[256:129], zll_main_multiply1749_inR49[128:1], zll_main_multiply1749_outR49);
  assign zll_main_multiply335_in = {zll_main_multiply389_in[255:128], zll_main_multiply389_in[127:0], (zll_main_multiply1749_inR49[0] == 1'h1) ? zll_main_multiply1749_outR49 : zll_main_multiply1792_outR111};
  assign id_inR335 = zll_main_multiply335_in[255:128];
  assign rewire_prelude_not_inR111 = id_inR335[0];
  ReWire_Prelude_not  instR446 (rewire_prelude_not_inR111[0], rewire_prelude_not_outR111);
  assign zll_main_multiply1785_inR111 = {zll_main_multiply335_in[255:128], rewire_prelude_not_outR111};
  ZLL_Main_multiply1785  instR447 (zll_main_multiply1785_inR111[128:1], zll_main_multiply1785_inR111[0], zll_main_multiply1785_outR111);
  assign zll_main_multiply295_in = {zll_main_multiply335_in[127:0], zll_main_multiply335_in[383:256], zll_main_multiply1785_outR111};
  assign id_inR336 = zll_main_multiply295_in[255:128];
  assign zll_main_multiply563_in = {zll_main_multiply295_in[383:256], zll_main_multiply295_in[255:128], zll_main_multiply295_in[127:0], id_inR336[15]};
  assign id_inR337 = zll_main_multiply563_in[256:129];
  assign zll_main_multiply1792_inR112 = {zll_main_multiply563_in[384:257], id_inR337[15]};
  ZLL_Main_multiply1792  instR448 (zll_main_multiply1792_inR112[128:1], zll_main_multiply1792_inR112[0], zll_main_multiply1792_outR112);
  assign zll_main_multiply1749_inR50 = {zll_main_multiply563_in[384:257], zll_main_multiply563_in[128:1], zll_main_multiply563_in[0]};
  ZLL_Main_multiply1749  instR449 (zll_main_multiply1749_inR50[256:129], zll_main_multiply1749_inR50[128:1], zll_main_multiply1749_outR50);
  assign zll_main_multiply1696_in = {zll_main_multiply295_in[255:128], zll_main_multiply295_in[127:0], (zll_main_multiply1749_inR50[0] == 1'h1) ? zll_main_multiply1749_outR50 : zll_main_multiply1792_outR112};
  assign id_inR338 = zll_main_multiply1696_in[255:128];
  assign rewire_prelude_not_inR112 = id_inR338[0];
  ReWire_Prelude_not  instR450 (rewire_prelude_not_inR112[0], rewire_prelude_not_outR112);
  assign zll_main_multiply1785_inR112 = {zll_main_multiply1696_in[255:128], rewire_prelude_not_outR112};
  ZLL_Main_multiply1785  instR451 (zll_main_multiply1785_inR112[128:1], zll_main_multiply1785_inR112[0], zll_main_multiply1785_outR112);
  assign zll_main_multiply1154_in = {zll_main_multiply1696_in[383:256], zll_main_multiply1696_in[127:0], zll_main_multiply1785_outR112};
  assign id_inR339 = zll_main_multiply1154_in[383:256];
  assign zll_main_multiply1017_in = {zll_main_multiply1154_in[127:0], zll_main_multiply1154_in[383:256], zll_main_multiply1154_in[255:128], id_inR339[14]};
  assign id_inR340 = zll_main_multiply1017_in[256:129];
  assign zll_main_multiply1792_inR113 = {zll_main_multiply1017_in[128:1], id_inR340[14]};
  ZLL_Main_multiply1792  instR452 (zll_main_multiply1792_inR113[128:1], zll_main_multiply1792_inR113[0], zll_main_multiply1792_outR113);
  assign zll_main_multiply1788_inR62 = {zll_main_multiply1017_in[384:257], zll_main_multiply1017_in[128:1], zll_main_multiply1017_in[0]};
  ZLL_Main_multiply1788  instR453 (zll_main_multiply1788_inR62[256:129], zll_main_multiply1788_inR62[128:1], zll_main_multiply1788_outR62);
  assign zll_main_multiply1568_in = {zll_main_multiply1154_in[127:0], zll_main_multiply1154_in[383:256], (zll_main_multiply1788_inR62[0] == 1'h1) ? zll_main_multiply1788_outR62 : zll_main_multiply1792_outR113};
  assign id_inR341 = zll_main_multiply1568_in[383:256];
  assign rewire_prelude_not_inR113 = id_inR341[0];
  ReWire_Prelude_not  instR454 (rewire_prelude_not_inR113[0], rewire_prelude_not_outR113);
  assign zll_main_multiply1785_inR113 = {zll_main_multiply1568_in[383:256], rewire_prelude_not_outR113};
  ZLL_Main_multiply1785  instR455 (zll_main_multiply1785_inR113[128:1], zll_main_multiply1785_inR113[0], zll_main_multiply1785_outR113);
  assign zll_main_multiply921_in = {zll_main_multiply1568_in[127:0], zll_main_multiply1568_in[255:128], zll_main_multiply1785_outR113};
  assign id_inR342 = zll_main_multiply921_in[255:128];
  assign zll_main_multiply576_in = {zll_main_multiply921_in[383:256], zll_main_multiply921_in[255:128], zll_main_multiply921_in[127:0], id_inR342[13]};
  assign id_inR343 = zll_main_multiply576_in[256:129];
  assign zll_main_multiply1792_inR114 = {zll_main_multiply576_in[384:257], id_inR343[13]};
  ZLL_Main_multiply1792  instR456 (zll_main_multiply1792_inR114[128:1], zll_main_multiply1792_inR114[0], zll_main_multiply1792_outR114);
  assign zll_main_multiply1749_inR51 = {zll_main_multiply576_in[384:257], zll_main_multiply576_in[128:1], zll_main_multiply576_in[0]};
  ZLL_Main_multiply1749  instR457 (zll_main_multiply1749_inR51[256:129], zll_main_multiply1749_inR51[128:1], zll_main_multiply1749_outR51);
  assign zll_main_multiply1358_in = {zll_main_multiply921_in[255:128], zll_main_multiply921_in[127:0], (zll_main_multiply1749_inR51[0] == 1'h1) ? zll_main_multiply1749_outR51 : zll_main_multiply1792_outR114};
  assign id_inR344 = zll_main_multiply1358_in[255:128];
  assign rewire_prelude_not_inR114 = id_inR344[0];
  ReWire_Prelude_not  instR458 (rewire_prelude_not_inR114[0], rewire_prelude_not_outR114);
  assign zll_main_multiply1785_inR114 = {zll_main_multiply1358_in[255:128], rewire_prelude_not_outR114};
  ZLL_Main_multiply1785  instR459 (zll_main_multiply1785_inR114[128:1], zll_main_multiply1785_inR114[0], zll_main_multiply1785_outR114);
  assign zll_main_multiply606_in = {zll_main_multiply1358_in[127:0], zll_main_multiply1358_in[383:256], zll_main_multiply1785_outR114};
  assign id_inR345 = zll_main_multiply606_in[255:128];
  assign zll_main_multiply567_in = {zll_main_multiply606_in[383:256], zll_main_multiply606_in[255:128], zll_main_multiply606_in[127:0], id_inR345[12]};
  assign id_inR346 = zll_main_multiply567_in[256:129];
  assign zll_main_multiply1792_inR115 = {zll_main_multiply567_in[384:257], id_inR346[12]};
  ZLL_Main_multiply1792  instR460 (zll_main_multiply1792_inR115[128:1], zll_main_multiply1792_inR115[0], zll_main_multiply1792_outR115);
  assign zll_main_multiply1749_inR52 = {zll_main_multiply567_in[384:257], zll_main_multiply567_in[128:1], zll_main_multiply567_in[0]};
  ZLL_Main_multiply1749  instR461 (zll_main_multiply1749_inR52[256:129], zll_main_multiply1749_inR52[128:1], zll_main_multiply1749_outR52);
  assign zll_main_multiply793_in = {zll_main_multiply606_in[255:128], zll_main_multiply606_in[127:0], (zll_main_multiply1749_inR52[0] == 1'h1) ? zll_main_multiply1749_outR52 : zll_main_multiply1792_outR115};
  assign id_inR347 = zll_main_multiply793_in[255:128];
  assign rewire_prelude_not_inR115 = id_inR347[0];
  ReWire_Prelude_not  instR462 (rewire_prelude_not_inR115[0], rewire_prelude_not_outR115);
  assign zll_main_multiply1785_inR115 = {zll_main_multiply793_in[255:128], rewire_prelude_not_outR115};
  ZLL_Main_multiply1785  instR463 (zll_main_multiply1785_inR115[128:1], zll_main_multiply1785_inR115[0], zll_main_multiply1785_outR115);
  assign zll_main_multiply636_in = {zll_main_multiply793_in[127:0], zll_main_multiply793_in[383:256], zll_main_multiply1785_outR115};
  assign id_inR348 = zll_main_multiply636_in[255:128];
  assign zll_main_multiply299_in = {zll_main_multiply636_in[127:0], zll_main_multiply636_in[383:256], zll_main_multiply636_in[255:128], id_inR348[11]};
  assign id_inR349 = zll_main_multiply299_in[128:1];
  assign zll_main_multiply1792_inR116 = {zll_main_multiply299_in[256:129], id_inR349[11]};
  ZLL_Main_multiply1792  instR464 (zll_main_multiply1792_inR116[128:1], zll_main_multiply1792_inR116[0], zll_main_multiply1792_outR116);
  assign zll_main_multiply1788_inR63 = {zll_main_multiply299_in[384:257], zll_main_multiply299_in[256:129], zll_main_multiply299_in[0]};
  ZLL_Main_multiply1788  instR465 (zll_main_multiply1788_inR63[256:129], zll_main_multiply1788_inR63[128:1], zll_main_multiply1788_outR63);
  assign zll_main_multiply1705_in = {zll_main_multiply636_in[127:0], zll_main_multiply636_in[255:128], (zll_main_multiply1788_inR63[0] == 1'h1) ? zll_main_multiply1788_outR63 : zll_main_multiply1792_outR116};
  assign id_inR350 = zll_main_multiply1705_in[383:256];
  assign rewire_prelude_not_inR116 = id_inR350[0];
  ReWire_Prelude_not  instR466 (rewire_prelude_not_inR116[0], rewire_prelude_not_outR116);
  assign zll_main_multiply1785_inR116 = {zll_main_multiply1705_in[383:256], rewire_prelude_not_outR116};
  ZLL_Main_multiply1785  instR467 (zll_main_multiply1785_inR116[128:1], zll_main_multiply1785_inR116[0], zll_main_multiply1785_outR116);
  assign zll_main_multiply439_in = {zll_main_multiply1705_in[127:0], zll_main_multiply1705_in[255:128], zll_main_multiply1785_outR116};
  assign id_inR351 = zll_main_multiply439_in[255:128];
  assign zll_main_multiply263_in = {zll_main_multiply439_in[127:0], zll_main_multiply439_in[383:256], zll_main_multiply439_in[255:128], id_inR351[10]};
  assign id_inR352 = zll_main_multiply263_in[128:1];
  assign zll_main_multiply1792_inR117 = {zll_main_multiply263_in[256:129], id_inR352[10]};
  ZLL_Main_multiply1792  instR468 (zll_main_multiply1792_inR117[128:1], zll_main_multiply1792_inR117[0], zll_main_multiply1792_outR117);
  assign zll_main_multiply1788_inR64 = {zll_main_multiply263_in[384:257], zll_main_multiply263_in[256:129], zll_main_multiply263_in[0]};
  ZLL_Main_multiply1788  instR469 (zll_main_multiply1788_inR64[256:129], zll_main_multiply1788_inR64[128:1], zll_main_multiply1788_outR64);
  assign zll_main_multiply1220_in = {zll_main_multiply439_in[127:0], zll_main_multiply439_in[255:128], (zll_main_multiply1788_inR64[0] == 1'h1) ? zll_main_multiply1788_outR64 : zll_main_multiply1792_outR117};
  assign id_inR353 = zll_main_multiply1220_in[383:256];
  assign rewire_prelude_not_inR117 = id_inR353[0];
  ReWire_Prelude_not  instR470 (rewire_prelude_not_inR117[0], rewire_prelude_not_outR117);
  assign zll_main_multiply1785_inR117 = {zll_main_multiply1220_in[383:256], rewire_prelude_not_outR117};
  ZLL_Main_multiply1785  instR471 (zll_main_multiply1785_inR117[128:1], zll_main_multiply1785_inR117[0], zll_main_multiply1785_outR117);
  assign zll_main_multiply430_in = {zll_main_multiply1220_in[127:0], zll_main_multiply1220_in[255:128], zll_main_multiply1785_outR117};
  assign id_inR354 = zll_main_multiply430_in[255:128];
  assign zll_main_multiply930_in = {zll_main_multiply430_in[383:256], zll_main_multiply430_in[255:128], zll_main_multiply430_in[127:0], id_inR354[9]};
  assign id_inR355 = zll_main_multiply930_in[256:129];
  assign zll_main_multiply1792_inR118 = {zll_main_multiply930_in[384:257], id_inR355[9]};
  ZLL_Main_multiply1792  instR472 (zll_main_multiply1792_inR118[128:1], zll_main_multiply1792_inR118[0], zll_main_multiply1792_outR118);
  assign zll_main_multiply1749_inR53 = {zll_main_multiply930_in[384:257], zll_main_multiply930_in[128:1], zll_main_multiply930_in[0]};
  ZLL_Main_multiply1749  instR473 (zll_main_multiply1749_inR53[256:129], zll_main_multiply1749_inR53[128:1], zll_main_multiply1749_outR53);
  assign zll_main_multiply443_in = {zll_main_multiply430_in[255:128], zll_main_multiply430_in[127:0], (zll_main_multiply1749_inR53[0] == 1'h1) ? zll_main_multiply1749_outR53 : zll_main_multiply1792_outR118};
  assign id_inR356 = zll_main_multiply443_in[255:128];
  assign rewire_prelude_not_inR118 = id_inR356[0];
  ReWire_Prelude_not  instR474 (rewire_prelude_not_inR118[0], rewire_prelude_not_outR118);
  assign zll_main_multiply1785_inR118 = {zll_main_multiply443_in[255:128], rewire_prelude_not_outR118};
  ZLL_Main_multiply1785  instR475 (zll_main_multiply1785_inR118[128:1], zll_main_multiply1785_inR118[0], zll_main_multiply1785_outR118);
  assign zll_main_multiply515_in = {zll_main_multiply443_in[127:0], zll_main_multiply443_in[383:256], zll_main_multiply1785_outR118};
  assign id_inR357 = zll_main_multiply515_in[255:128];
  assign zll_main_multiply763_in = {zll_main_multiply515_in[383:256], zll_main_multiply515_in[127:0], zll_main_multiply515_in[255:128], id_inR357[8]};
  assign id_inR358 = zll_main_multiply763_in[128:1];
  assign zll_main_multiply1792_inR119 = {zll_main_multiply763_in[384:257], id_inR358[8]};
  ZLL_Main_multiply1792  instR476 (zll_main_multiply1792_inR119[128:1], zll_main_multiply1792_inR119[0], zll_main_multiply1792_outR119);
  assign zll_main_multiply1749_inR54 = {zll_main_multiply763_in[384:257], zll_main_multiply763_in[256:129], zll_main_multiply763_in[0]};
  ZLL_Main_multiply1749  instR477 (zll_main_multiply1749_inR54[256:129], zll_main_multiply1749_inR54[128:1], zll_main_multiply1749_outR54);
  assign zll_main_multiply1725_in = {zll_main_multiply515_in[127:0], zll_main_multiply515_in[255:128], (zll_main_multiply1749_inR54[0] == 1'h1) ? zll_main_multiply1749_outR54 : zll_main_multiply1792_outR119};
  assign id_inR359 = zll_main_multiply1725_in[383:256];
  assign rewire_prelude_not_inR119 = id_inR359[0];
  ReWire_Prelude_not  instR478 (rewire_prelude_not_inR119[0], rewire_prelude_not_outR119);
  assign zll_main_multiply1785_inR119 = {zll_main_multiply1725_in[383:256], rewire_prelude_not_outR119};
  ZLL_Main_multiply1785  instR479 (zll_main_multiply1785_inR119[128:1], zll_main_multiply1785_inR119[0], zll_main_multiply1785_outR119);
  assign zll_main_multiply1425_in = {zll_main_multiply1725_in[127:0], zll_main_multiply1725_in[255:128], zll_main_multiply1785_outR119};
  assign id_inR360 = zll_main_multiply1425_in[255:128];
  assign zll_main_multiply1784_in = {zll_main_multiply1425_in[383:256], zll_main_multiply1425_in[255:128], zll_main_multiply1425_in[127:0], id_inR360[7]};
  assign id_inR361 = zll_main_multiply1784_in[256:129];
  assign zll_main_multiply1792_inR120 = {zll_main_multiply1784_in[384:257], id_inR361[7]};
  ZLL_Main_multiply1792  instR480 (zll_main_multiply1792_inR120[128:1], zll_main_multiply1792_inR120[0], zll_main_multiply1792_outR120);
  assign zll_main_multiply1749_inR55 = {zll_main_multiply1784_in[384:257], zll_main_multiply1784_in[128:1], zll_main_multiply1784_in[0]};
  ZLL_Main_multiply1749  instR481 (zll_main_multiply1749_inR55[256:129], zll_main_multiply1749_inR55[128:1], zll_main_multiply1749_outR55);
  assign zll_main_multiply1306_in = {zll_main_multiply1425_in[255:128], zll_main_multiply1425_in[127:0], (zll_main_multiply1749_inR55[0] == 1'h1) ? zll_main_multiply1749_outR55 : zll_main_multiply1792_outR120};
  assign id_inR362 = zll_main_multiply1306_in[255:128];
  assign rewire_prelude_not_inR120 = id_inR362[0];
  ReWire_Prelude_not  instR482 (rewire_prelude_not_inR120[0], rewire_prelude_not_outR120);
  assign zll_main_multiply1785_inR120 = {zll_main_multiply1306_in[255:128], rewire_prelude_not_outR120};
  ZLL_Main_multiply1785  instR483 (zll_main_multiply1785_inR120[128:1], zll_main_multiply1785_inR120[0], zll_main_multiply1785_outR120);
  assign zll_main_multiply1407_in = {zll_main_multiply1306_in[127:0], zll_main_multiply1306_in[383:256], zll_main_multiply1785_outR120};
  assign id_inR363 = zll_main_multiply1407_in[255:128];
  assign zll_main_multiply692_in = {zll_main_multiply1407_in[127:0], zll_main_multiply1407_in[383:256], zll_main_multiply1407_in[255:128], id_inR363[6]};
  assign id_inR364 = zll_main_multiply692_in[128:1];
  assign zll_main_multiply1792_inR121 = {zll_main_multiply692_in[256:129], id_inR364[6]};
  ZLL_Main_multiply1792  instR484 (zll_main_multiply1792_inR121[128:1], zll_main_multiply1792_inR121[0], zll_main_multiply1792_outR121);
  assign zll_main_multiply1788_inR65 = {zll_main_multiply692_in[384:257], zll_main_multiply692_in[256:129], zll_main_multiply692_in[0]};
  ZLL_Main_multiply1788  instR485 (zll_main_multiply1788_inR65[256:129], zll_main_multiply1788_inR65[128:1], zll_main_multiply1788_outR65);
  assign zll_main_multiply850_in = {zll_main_multiply1407_in[127:0], zll_main_multiply1407_in[255:128], (zll_main_multiply1788_inR65[0] == 1'h1) ? zll_main_multiply1788_outR65 : zll_main_multiply1792_outR121};
  assign id_inR365 = zll_main_multiply850_in[383:256];
  assign rewire_prelude_not_inR121 = id_inR365[0];
  ReWire_Prelude_not  instR486 (rewire_prelude_not_inR121[0], rewire_prelude_not_outR121);
  assign zll_main_multiply1785_inR121 = {zll_main_multiply850_in[383:256], rewire_prelude_not_outR121};
  ZLL_Main_multiply1785  instR487 (zll_main_multiply1785_inR121[128:1], zll_main_multiply1785_inR121[0], zll_main_multiply1785_outR121);
  assign zll_main_multiply392_in = {zll_main_multiply850_in[255:128], zll_main_multiply850_in[127:0], zll_main_multiply1785_outR121};
  assign id_inR366 = zll_main_multiply392_in[383:256];
  assign zll_main_multiply887_in = {zll_main_multiply392_in[127:0], zll_main_multiply392_in[383:256], zll_main_multiply392_in[255:128], id_inR366[5]};
  assign id_inR367 = zll_main_multiply887_in[256:129];
  assign zll_main_multiply1792_inR122 = {zll_main_multiply887_in[128:1], id_inR367[5]};
  ZLL_Main_multiply1792  instR488 (zll_main_multiply1792_inR122[128:1], zll_main_multiply1792_inR122[0], zll_main_multiply1792_outR122);
  assign zll_main_multiply1788_inR66 = {zll_main_multiply887_in[384:257], zll_main_multiply887_in[128:1], zll_main_multiply887_in[0]};
  ZLL_Main_multiply1788  instR489 (zll_main_multiply1788_inR66[256:129], zll_main_multiply1788_inR66[128:1], zll_main_multiply1788_outR66);
  assign zll_main_multiply1426_in = {zll_main_multiply392_in[127:0], zll_main_multiply392_in[383:256], (zll_main_multiply1788_inR66[0] == 1'h1) ? zll_main_multiply1788_outR66 : zll_main_multiply1792_outR122};
  assign id_inR368 = zll_main_multiply1426_in[383:256];
  assign rewire_prelude_not_inR122 = id_inR368[0];
  ReWire_Prelude_not  instR490 (rewire_prelude_not_inR122[0], rewire_prelude_not_outR122);
  assign zll_main_multiply1785_inR122 = {zll_main_multiply1426_in[383:256], rewire_prelude_not_outR122};
  ZLL_Main_multiply1785  instR491 (zll_main_multiply1785_inR122[128:1], zll_main_multiply1785_inR122[0], zll_main_multiply1785_outR122);
  assign zll_main_multiply1704_in = {zll_main_multiply1426_in[127:0], zll_main_multiply1426_in[255:128], zll_main_multiply1785_outR122};
  assign id_inR369 = zll_main_multiply1704_in[255:128];
  assign zll_main_multiply758_in = {zll_main_multiply1704_in[383:256], zll_main_multiply1704_in[127:0], zll_main_multiply1704_in[255:128], id_inR369[4]};
  assign id_inR370 = zll_main_multiply758_in[128:1];
  assign zll_main_multiply1792_inR123 = {zll_main_multiply758_in[384:257], id_inR370[4]};
  ZLL_Main_multiply1792  instR492 (zll_main_multiply1792_inR123[128:1], zll_main_multiply1792_inR123[0], zll_main_multiply1792_outR123);
  assign zll_main_multiply1749_inR56 = {zll_main_multiply758_in[384:257], zll_main_multiply758_in[256:129], zll_main_multiply758_in[0]};
  ZLL_Main_multiply1749  instR493 (zll_main_multiply1749_inR56[256:129], zll_main_multiply1749_inR56[128:1], zll_main_multiply1749_outR56);
  assign zll_main_multiply537_in = {zll_main_multiply1704_in[127:0], zll_main_multiply1704_in[255:128], (zll_main_multiply1749_inR56[0] == 1'h1) ? zll_main_multiply1749_outR56 : zll_main_multiply1792_outR123};
  assign id_inR371 = zll_main_multiply537_in[383:256];
  assign rewire_prelude_not_inR123 = id_inR371[0];
  ReWire_Prelude_not  instR494 (rewire_prelude_not_inR123[0], rewire_prelude_not_outR123);
  assign zll_main_multiply1785_inR123 = {zll_main_multiply537_in[383:256], rewire_prelude_not_outR123};
  ZLL_Main_multiply1785  instR495 (zll_main_multiply1785_inR123[128:1], zll_main_multiply1785_inR123[0], zll_main_multiply1785_outR123);
  assign zll_main_multiply446_in = {zll_main_multiply537_in[255:128], zll_main_multiply537_in[127:0], zll_main_multiply1785_outR123};
  assign id_inR372 = zll_main_multiply446_in[383:256];
  assign zll_main_multiply1681_in = {zll_main_multiply446_in[127:0], zll_main_multiply446_in[383:256], zll_main_multiply446_in[255:128], id_inR372[3]};
  assign id_inR373 = zll_main_multiply1681_in[256:129];
  assign zll_main_multiply1792_inR124 = {zll_main_multiply1681_in[128:1], id_inR373[3]};
  ZLL_Main_multiply1792  instR496 (zll_main_multiply1792_inR124[128:1], zll_main_multiply1792_inR124[0], zll_main_multiply1792_outR124);
  assign zll_main_multiply1788_inR67 = {zll_main_multiply1681_in[384:257], zll_main_multiply1681_in[128:1], zll_main_multiply1681_in[0]};
  ZLL_Main_multiply1788  instR497 (zll_main_multiply1788_inR67[256:129], zll_main_multiply1788_inR67[128:1], zll_main_multiply1788_outR67);
  assign zll_main_multiply1125_in = {zll_main_multiply446_in[127:0], zll_main_multiply446_in[383:256], (zll_main_multiply1788_inR67[0] == 1'h1) ? zll_main_multiply1788_outR67 : zll_main_multiply1792_outR124};
  assign id_inR374 = zll_main_multiply1125_in[383:256];
  assign rewire_prelude_not_inR124 = id_inR374[0];
  ReWire_Prelude_not  instR498 (rewire_prelude_not_inR124[0], rewire_prelude_not_outR124);
  assign zll_main_multiply1785_inR124 = {zll_main_multiply1125_in[383:256], rewire_prelude_not_outR124};
  ZLL_Main_multiply1785  instR499 (zll_main_multiply1785_inR124[128:1], zll_main_multiply1785_inR124[0], zll_main_multiply1785_outR124);
  assign zll_main_multiply1429_in = {zll_main_multiply1125_in[127:0], zll_main_multiply1125_in[255:128], zll_main_multiply1785_outR124};
  assign id_inR375 = zll_main_multiply1429_in[255:128];
  assign zll_main_multiply881_in = {zll_main_multiply1429_in[383:256], zll_main_multiply1429_in[255:128], zll_main_multiply1429_in[127:0], id_inR375[2]};
  assign id_inR376 = zll_main_multiply881_in[256:129];
  assign zll_main_multiply1792_inR125 = {zll_main_multiply881_in[384:257], id_inR376[2]};
  ZLL_Main_multiply1792  instR500 (zll_main_multiply1792_inR125[128:1], zll_main_multiply1792_inR125[0], zll_main_multiply1792_outR125);
  assign zll_main_multiply1749_inR57 = {zll_main_multiply881_in[384:257], zll_main_multiply881_in[128:1], zll_main_multiply881_in[0]};
  ZLL_Main_multiply1749  instR501 (zll_main_multiply1749_inR57[256:129], zll_main_multiply1749_inR57[128:1], zll_main_multiply1749_outR57);
  assign zll_main_multiply1113_in = {zll_main_multiply1429_in[255:128], zll_main_multiply1429_in[127:0], (zll_main_multiply1749_inR57[0] == 1'h1) ? zll_main_multiply1749_outR57 : zll_main_multiply1792_outR125};
  assign id_inR377 = zll_main_multiply1113_in[255:128];
  assign rewire_prelude_not_inR125 = id_inR377[0];
  ReWire_Prelude_not  instR502 (rewire_prelude_not_inR125[0], rewire_prelude_not_outR125);
  assign zll_main_multiply1785_inR125 = {zll_main_multiply1113_in[255:128], rewire_prelude_not_outR125};
  ZLL_Main_multiply1785  instR503 (zll_main_multiply1785_inR125[128:1], zll_main_multiply1785_inR125[0], zll_main_multiply1785_outR125);
  assign zll_main_multiply1192_in = {zll_main_multiply1113_in[383:256], zll_main_multiply1113_in[127:0], zll_main_multiply1785_outR125};
  assign id_inR378 = zll_main_multiply1192_in[383:256];
  assign zll_main_multiply695_in = {zll_main_multiply1192_in[127:0], zll_main_multiply1192_in[383:256], zll_main_multiply1192_in[255:128], id_inR378[1]};
  assign id_inR379 = zll_main_multiply695_in[256:129];
  assign zll_main_multiply1792_inR126 = {zll_main_multiply695_in[128:1], id_inR379[1]};
  ZLL_Main_multiply1792  instR504 (zll_main_multiply1792_inR126[128:1], zll_main_multiply1792_inR126[0], zll_main_multiply1792_outR126);
  assign zll_main_multiply1788_inR68 = {zll_main_multiply695_in[384:257], zll_main_multiply695_in[128:1], zll_main_multiply695_in[0]};
  ZLL_Main_multiply1788  instR505 (zll_main_multiply1788_inR68[256:129], zll_main_multiply1788_inR68[128:1], zll_main_multiply1788_outR68);
  assign zll_main_multiply360_in = {zll_main_multiply1192_in[127:0], zll_main_multiply1192_in[383:256], (zll_main_multiply1788_inR68[0] == 1'h1) ? zll_main_multiply1788_outR68 : zll_main_multiply1792_outR126};
  assign id_inR380 = zll_main_multiply360_in[383:256];
  assign rewire_prelude_not_inR126 = id_inR380[0];
  ReWire_Prelude_not  instR506 (rewire_prelude_not_inR126[0], rewire_prelude_not_outR126);
  assign zll_main_multiply1785_inR126 = {zll_main_multiply360_in[383:256], rewire_prelude_not_outR126};
  ZLL_Main_multiply1785  instR507 (zll_main_multiply1785_inR126[128:1], zll_main_multiply1785_inR126[0], zll_main_multiply1785_outR126);
  assign zll_main_multiply767_in = {zll_main_multiply360_in[127:0], zll_main_multiply360_in[255:128], zll_main_multiply1785_outR126};
  assign id_inR381 = zll_main_multiply767_in[255:128];
  assign zll_main_multiply608_in = {zll_main_multiply767_in[127:0], zll_main_multiply767_in[383:256], zll_main_multiply767_in[255:128], id_inR381[0]};
  assign id_inR382 = zll_main_multiply608_in[128:1];
  assign zll_main_multiply1792_inR127 = {zll_main_multiply608_in[256:129], id_inR382[0]};
  ZLL_Main_multiply1792  instR508 (zll_main_multiply1792_inR127[128:1], zll_main_multiply1792_inR127[0], zll_main_multiply1792_outR127);
  assign zll_main_multiply1788_inR69 = {zll_main_multiply608_in[384:257], zll_main_multiply608_in[256:129], zll_main_multiply608_in[0]};
  ZLL_Main_multiply1788  instR509 (zll_main_multiply1788_inR69[256:129], zll_main_multiply1788_inR69[128:1], zll_main_multiply1788_outR69);
  assign {__continue, __out0} = (zll_main_multiply1788_inR69[0] == 1'h1) ? zll_main_multiply1788_outR69 : zll_main_multiply1792_outR127;
endmodule

module ZLL_Main_multiply1792 (input logic [127:0] arg0,
  input logic [0:0] arg1,
  output logic [127:0] res);
  logic [128:0] id_in;
  assign id_in = {arg0, arg1};
  assign res = id_in[128:1];
endmodule

module ZLL_Main_multiply1788 (input logic [127:0] arg0,
  input logic [127:0] arg1,
  output logic [127:0] res);
  logic [255:0] binop_in;
  assign binop_in = {arg1, arg0};
  assign res = binop_in[255:128] ^ binop_in[127:0];
endmodule

module ZLL_Main_multiply1785 (input logic [127:0] arg0,
  input logic [0:0] arg1,
  output logic [127:0] res);
  logic [127:0] id_in;
  logic [0:0] rewire_prelude_not_in;
  logic [0:0] rewire_prelude_not_out;
  logic [128:0] zll_main_multiply1780_in;
  logic [128:0] zll_main_multiply1767_in;
  logic [255:0] binop_in;
  logic [255:0] binop_inR1;
  logic [128:0] zll_main_multiply1779_in;
  logic [255:0] binop_inR2;
  assign id_in = arg0;
  assign rewire_prelude_not_in = id_in[0];
  ReWire_Prelude_not  inst (rewire_prelude_not_in[0], rewire_prelude_not_out);
  assign zll_main_multiply1780_in = {arg0, rewire_prelude_not_out};
  assign zll_main_multiply1767_in = {zll_main_multiply1780_in[128:1], zll_main_multiply1780_in[0]};
  assign binop_in = {zll_main_multiply1767_in[128:1], 128'h1};
  assign binop_inR1 = {binop_in[255:128] >> binop_in[127:0], {8'he1, {7'h78{1'h0}}}};
  assign zll_main_multiply1779_in = {arg0, arg1};
  assign binop_inR2 = {zll_main_multiply1779_in[128:1], 128'h1};
  assign res = (zll_main_multiply1779_in[0] == 1'h1) ? (binop_inR2[255:128] >> binop_inR2[127:0]) : (binop_inR1[255:128] ^ binop_inR1[127:0]);
endmodule

module ZLL_Main_multiply1749 (input logic [127:0] arg0,
  input logic [127:0] arg1,
  output logic [127:0] res);
  logic [255:0] binop_in;
  assign binop_in = {arg0, arg1};
  assign res = binop_in[255:128] ^ binop_in[127:0];
endmodule

module ReWire_Prelude_not (input logic [0:0] arg0,
  output logic [0:0] res);
  logic [1:0] zll_rewire_prelude_not_in;
  logic [0:0] lit_in;
  assign zll_rewire_prelude_not_in = {arg0, arg0};
  assign lit_in = zll_rewire_prelude_not_in[0];
  assign res = (lit_in[0] == 1'h1) ? 1'h0 : 1'h1;
endmodule