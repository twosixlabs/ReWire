module top_level (input logic [6:0] __in0,
  output logic [4:0] __out0);
  logic [6:0] zll_main_loop1_in;
  logic [6:0] zll_main_compute1_in;
  logic [6:0] resize_in;
  logic [6:0] resize_inR1;
  logic [255:0] binop_in;
  logic [127:0] resize_inR2;
  logic [4:0] zll_main_compute2_in;
  logic [9:0] zll_main_compute4_in;
  logic [9:0] zll_main_compute6_in;
  logic [9:0] zll_main_compute_in;
  logic [4:0] resize_inR3;
  logic [4:0] resize_inR4;
  logic [255:0] binop_inR1;
  logic [255:0] binop_inR2;
  logic [127:0] resize_inR5;
  logic [5:0] zll_main_loop2_in;
  logic [5:0] zll_main_loop3_in;
  logic [0:0] __continue;
  assign zll_main_loop1_in = __in0;
  assign zll_main_compute1_in = zll_main_loop1_in[6:0];
  assign resize_in = zll_main_compute1_in[6:0];
  assign resize_inR1 = resize_in[6:0];
  assign binop_in = {128'(resize_inR1[6:0]), 128'h14};
  assign resize_inR2 = binop_in[255:128] % binop_in[127:0];
  assign zll_main_compute2_in = resize_inR2[4:0];
  assign zll_main_compute4_in = {zll_main_compute2_in[4:0], 5'h6};
  assign zll_main_compute6_in = {zll_main_compute4_in[9:5], zll_main_compute4_in[4:0]};
  assign zll_main_compute_in = zll_main_compute6_in[9:0];
  assign resize_inR3 = zll_main_compute_in[9:5];
  assign resize_inR4 = zll_main_compute_in[4:0];
  assign binop_inR1 = {128'(resize_inR3[4:0]), 128'(resize_inR4[4:0])};
  assign binop_inR2 = {binop_inR1[255:128] + binop_inR1[127:0], 128'h14};
  assign resize_inR5 = binop_inR2[255:128] % binop_inR2[127:0];
  assign zll_main_loop2_in = {1'h0, resize_inR5[4:0]};
  assign zll_main_loop3_in = zll_main_loop2_in[5:0];
  assign {__continue, __out0} = {1'h1, zll_main_loop3_in[4:0]};
endmodule