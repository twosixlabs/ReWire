module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [63:0] __in0,
  input logic [63:0] __in1,
  output logic [63:0] __out0,
  output logic [63:0] __out1);
  logic [128:0] gzdLLzicase16315;
  logic [129:0] callRes;
  logic [128:0] gzdLLzicase16315R1;
  logic [129:0] callResR1;
  logic [0:0] __continue;
  logic [0:0] __resumption_tag;
  logic [0:0] __resumption_tag_next;
  assign gzdLLzicase16315 = {__resumption_tag, {__in0, __in1}};
  zdLLzicase16315  zdLLzicase16315 (gzdLLzicase16315[127:0], callRes);
  assign gzdLLzicase16315R1 = {__resumption_tag, {__in0, __in1}};
  zdLLzicase16315  zdLLzicase16315R1 (gzdLLzicase16315R1[127:0], callResR1);
  assign {__continue, __out0, __out1, __resumption_tag_next} = (gzdLLzicase16315R1[128] == 1'h0) ? callResR1 : callRes;
  initial __resumption_tag <= 1'h1;
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      __resumption_tag <= 1'h1;
    end else begin
      __resumption_tag <= __resumption_tag_next;
    end
  end
endmodule

module zdLLzicase16053 (input logic [63:0] arg0,
  input logic [2:0] arg1,
  output logic [7:0] res);
  logic [63:0] resizze;
  logic [2:0] resizzeR1;
  logic [255:0] binOp;
  logic [255:0] binOpR1;
  logic [127:0] resizzeR2;
  logic [2:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR6;
  logic [2:0] resizzeR7;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [127:0] resizzeR8;
  assign resizze = arg0;
  assign resizzeR1 = arg1;
  assign binOp = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign binOpR1 = {binOp[255:128] - binOp[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR2 = binOpR1[255:128] % binOpR1[127:0];
  assign resizzeR3 = resizzeR2[2:0];
  assign binOpR2 = {128'(resizzeR3[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR3 = {binOpR2[255:128] * binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[2:0];
  assign binOpR4 = {128'(resizzeR5[2:0]), 128'h00000000000000000000000000000001};
  assign binOpR5 = {binOpR4[255:128] + binOpR4[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR6 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR7 = resizzeR6[2:0];
  assign binOpR6 = {128'h00000000000000000000000000000008, 128'(resizzeR7[2:0])};
  assign binOpR7 = {binOpR6[255:128] - binOpR6[127:0], 128'h00000000000000000000000000000001};
  assign binOpR8 = {binOpR7[255:128] - binOpR7[127:0], 128'h00000000000000000000000000000008};
  assign binOpR9 = {128'(resizze[63:0]), binOpR8[255:128] * binOpR8[127:0]};
  assign resizzeR8 = binOpR9[255:128] >> binOpR9[127:0];
  assign res = resizzeR8[7:0];
endmodule

module zdLLzicase16056 (input logic [63:0] arg0,
  input logic [2:0] arg1,
  output logic [7:0] res);
  logic [63:0] resizze;
  logic [2:0] resizzeR1;
  logic [255:0] binOp;
  logic [255:0] binOpR1;
  logic [127:0] resizzeR2;
  logic [2:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [127:0] resizzeR6;
  assign resizze = arg0;
  assign resizzeR1 = arg1;
  assign binOp = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR1 = {binOp[255:128] * binOp[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR2 = binOpR1[255:128] % binOpR1[127:0];
  assign resizzeR3 = resizzeR2[2:0];
  assign binOpR2 = {128'(resizzeR3[2:0]), 128'h00000000000000000000000000000001};
  assign binOpR3 = {binOpR2[255:128] + binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[2:0];
  assign binOpR4 = {128'h00000000000000000000000000000008, 128'(resizzeR5[2:0])};
  assign binOpR5 = {binOpR4[255:128] - binOpR4[127:0], 128'h00000000000000000000000000000001};
  assign binOpR6 = {binOpR5[255:128] - binOpR5[127:0], 128'h00000000000000000000000000000008};
  assign binOpR7 = {128'(resizze[63:0]), binOpR6[255:128] * binOpR6[127:0]};
  assign resizzeR6 = binOpR7[255:128] >> binOpR7[127:0];
  assign res = resizzeR6[7:0];
endmodule

module zdLLzicase16063 (input logic [63:0] arg0,
  input logic [2:0] arg1,
  output logic [7:0] res);
  logic [63:0] resizze;
  logic [2:0] resizzeR1;
  logic [255:0] binOp;
  logic [255:0] binOpR1;
  logic [127:0] resizzeR2;
  logic [2:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [127:0] resizzeR6;
  assign resizze = arg0;
  assign resizzeR1 = arg1;
  assign binOp = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign binOpR1 = {binOp[255:128] - binOp[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR2 = binOpR1[255:128] % binOpR1[127:0];
  assign resizzeR3 = resizzeR2[2:0];
  assign binOpR2 = {128'(resizzeR3[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR3 = {binOpR2[255:128] * binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[2:0];
  assign binOpR4 = {128'h00000000000000000000000000000008, 128'(resizzeR5[2:0])};
  assign binOpR5 = {binOpR4[255:128] - binOpR4[127:0], 128'h00000000000000000000000000000001};
  assign binOpR6 = {binOpR5[255:128] - binOpR5[127:0], 128'h00000000000000000000000000000008};
  assign binOpR7 = {128'(resizze[63:0]), binOpR6[255:128] * binOpR6[127:0]};
  assign resizzeR6 = binOpR7[255:128] >> binOpR7[127:0];
  assign res = resizzeR6[7:0];
endmodule

module zdLLzicase16066 (input logic [63:0] arg0,
  input logic [2:0] arg1,
  output logic [7:0] res);
  logic [63:0] resizze;
  logic [2:0] resizzeR1;
  logic [255:0] binOp;
  logic [255:0] binOpR1;
  logic [127:0] resizzeR2;
  logic [2:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR4;
  assign resizze = arg0;
  assign resizzeR1 = arg1;
  assign binOp = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR1 = {binOp[255:128] * binOp[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR2 = binOpR1[255:128] % binOpR1[127:0];
  assign resizzeR3 = resizzeR2[2:0];
  assign binOpR2 = {128'h00000000000000000000000000000008, 128'(resizzeR3[2:0])};
  assign binOpR3 = {binOpR2[255:128] - binOpR2[127:0], 128'h00000000000000000000000000000001};
  assign binOpR4 = {binOpR3[255:128] - binOpR3[127:0], 128'h00000000000000000000000000000008};
  assign binOpR5 = {128'(resizze[63:0]), binOpR4[255:128] * binOpR4[127:0]};
  assign resizzeR4 = binOpR5[255:128] >> binOpR5[127:0];
  assign res = resizzeR4[7:0];
endmodule

module zdLLzicase16315 (input logic [127:0] arg0,
  output logic [129:0] res);
  logic [127:0] gMainziloop;
  logic [127:0] gMainzicompute;
  logic [127:0] gzdLLzicase16205;
  logic [130:0] gzdLLzilambda16126;
  logic [7:0] callRes;
  logic [130:0] gzdLLzilambda16126R1;
  logic [7:0] callResR1;
  logic [130:0] gzdLLzilambda16126R2;
  logic [7:0] callResR2;
  logic [130:0] gzdLLzilambda16126R3;
  logic [7:0] callResR3;
  logic [130:0] gzdLLzilambda16126R4;
  logic [7:0] callResR4;
  logic [130:0] gzdLLzilambda16126R5;
  logic [7:0] callResR5;
  logic [130:0] gzdLLzilambda16126R6;
  logic [7:0] callResR6;
  logic [130:0] gzdLLzilambda16126R7;
  logic [7:0] callResR7;
  logic [130:0] gzdLLzilambda16202;
  logic [7:0] callResR8;
  logic [130:0] gzdLLzilambda16202R1;
  logic [7:0] callResR9;
  logic [130:0] gzdLLzilambda16202R2;
  logic [7:0] callResR10;
  logic [130:0] gzdLLzilambda16202R3;
  logic [7:0] callResR11;
  logic [130:0] gzdLLzilambda16202R4;
  logic [7:0] callResR12;
  logic [130:0] gzdLLzilambda16202R5;
  logic [7:0] callResR13;
  logic [130:0] gzdLLzilambda16202R6;
  logic [7:0] callResR14;
  logic [130:0] gzdLLzilambda16202R7;
  logic [7:0] callResR15;
  logic [129:0] gzdLLzilambda16321;
  logic [129:0] gzdLLzicase16319;
  logic [127:0] gzdLLzilambda16209;
  assign gMainziloop = arg0;
  assign gMainzicompute = gMainziloop[127:0];
  assign gzdLLzicase16205 = gMainzicompute[127:0];
  assign gzdLLzilambda16126 = {gzdLLzicase16205[127:64], gzdLLzicase16205[63:0], 3'h0};
  zdLLzilambda16126  zdLLzilambda16126 (gzdLLzilambda16126[130:67], gzdLLzilambda16126[66:3], gzdLLzilambda16126[2:0], callRes);
  assign gzdLLzilambda16126R1 = {gzdLLzicase16205[127:64], gzdLLzicase16205[63:0], 3'h1};
  zdLLzilambda16126  zdLLzilambda16126R1 (gzdLLzilambda16126R1[130:67], gzdLLzilambda16126R1[66:3], gzdLLzilambda16126R1[2:0], callResR1);
  assign gzdLLzilambda16126R2 = {gzdLLzicase16205[127:64], gzdLLzicase16205[63:0], 3'h2};
  zdLLzilambda16126  zdLLzilambda16126R2 (gzdLLzilambda16126R2[130:67], gzdLLzilambda16126R2[66:3], gzdLLzilambda16126R2[2:0], callResR2);
  assign gzdLLzilambda16126R3 = {gzdLLzicase16205[127:64], gzdLLzicase16205[63:0], 3'h3};
  zdLLzilambda16126  zdLLzilambda16126R3 (gzdLLzilambda16126R3[130:67], gzdLLzilambda16126R3[66:3], gzdLLzilambda16126R3[2:0], callResR3);
  assign gzdLLzilambda16126R4 = {gzdLLzicase16205[127:64], gzdLLzicase16205[63:0], 3'h4};
  zdLLzilambda16126  zdLLzilambda16126R4 (gzdLLzilambda16126R4[130:67], gzdLLzilambda16126R4[66:3], gzdLLzilambda16126R4[2:0], callResR4);
  assign gzdLLzilambda16126R5 = {gzdLLzicase16205[127:64], gzdLLzicase16205[63:0], 3'h5};
  zdLLzilambda16126  zdLLzilambda16126R5 (gzdLLzilambda16126R5[130:67], gzdLLzilambda16126R5[66:3], gzdLLzilambda16126R5[2:0], callResR5);
  assign gzdLLzilambda16126R6 = {gzdLLzicase16205[127:64], gzdLLzicase16205[63:0], 3'h6};
  zdLLzilambda16126  zdLLzilambda16126R6 (gzdLLzilambda16126R6[130:67], gzdLLzilambda16126R6[66:3], gzdLLzilambda16126R6[2:0], callResR6);
  assign gzdLLzilambda16126R7 = {gzdLLzicase16205[127:64], gzdLLzicase16205[63:0], 3'h7};
  zdLLzilambda16126  zdLLzilambda16126R7 (gzdLLzilambda16126R7[130:67], gzdLLzilambda16126R7[66:3], gzdLLzilambda16126R7[2:0], callResR7);
  assign gzdLLzilambda16202 = {gzdLLzicase16205[127:64], gzdLLzicase16205[63:0], 3'h0};
  zdLLzilambda16202  zdLLzilambda16202 (gzdLLzilambda16202[130:67], gzdLLzilambda16202[66:3], gzdLLzilambda16202[2:0], callResR8);
  assign gzdLLzilambda16202R1 = {gzdLLzicase16205[127:64], gzdLLzicase16205[63:0], 3'h1};
  zdLLzilambda16202  zdLLzilambda16202R1 (gzdLLzilambda16202R1[130:67], gzdLLzilambda16202R1[66:3], gzdLLzilambda16202R1[2:0], callResR9);
  assign gzdLLzilambda16202R2 = {gzdLLzicase16205[127:64], gzdLLzicase16205[63:0], 3'h2};
  zdLLzilambda16202  zdLLzilambda16202R2 (gzdLLzilambda16202R2[130:67], gzdLLzilambda16202R2[66:3], gzdLLzilambda16202R2[2:0], callResR10);
  assign gzdLLzilambda16202R3 = {gzdLLzicase16205[127:64], gzdLLzicase16205[63:0], 3'h3};
  zdLLzilambda16202  zdLLzilambda16202R3 (gzdLLzilambda16202R3[130:67], gzdLLzilambda16202R3[66:3], gzdLLzilambda16202R3[2:0], callResR11);
  assign gzdLLzilambda16202R4 = {gzdLLzicase16205[127:64], gzdLLzicase16205[63:0], 3'h4};
  zdLLzilambda16202  zdLLzilambda16202R4 (gzdLLzilambda16202R4[130:67], gzdLLzilambda16202R4[66:3], gzdLLzilambda16202R4[2:0], callResR12);
  assign gzdLLzilambda16202R5 = {gzdLLzicase16205[127:64], gzdLLzicase16205[63:0], 3'h5};
  zdLLzilambda16202  zdLLzilambda16202R5 (gzdLLzilambda16202R5[130:67], gzdLLzilambda16202R5[66:3], gzdLLzilambda16202R5[2:0], callResR13);
  assign gzdLLzilambda16202R6 = {gzdLLzicase16205[127:64], gzdLLzicase16205[63:0], 3'h6};
  zdLLzilambda16202  zdLLzilambda16202R6 (gzdLLzilambda16202R6[130:67], gzdLLzilambda16202R6[66:3], gzdLLzilambda16202R6[2:0], callResR14);
  assign gzdLLzilambda16202R7 = {gzdLLzicase16205[127:64], gzdLLzicase16205[63:0], 3'h7};
  zdLLzilambda16202  zdLLzilambda16202R7 (gzdLLzilambda16202R7[130:67], gzdLLzilambda16202R7[66:3], gzdLLzilambda16202R7[2:0], callResR15);
  assign gzdLLzilambda16321 = {2'h0, {callRes, callResR1, callResR2, callResR3, callResR4, callResR5, callResR6, callResR7, callResR8, callResR9, callResR10, callResR11, callResR12, callResR13, callResR14, callResR15}};
  assign gzdLLzicase16319 = gzdLLzilambda16321[129:0];
  assign gzdLLzilambda16209 = gzdLLzicase16319[127:0];
  assign res = {1'h1, gzdLLzilambda16209[127:0], 1'h0};
endmodule

module zdLLzilambda16060 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [67:0] gzdLLzicase16053;
  logic [7:0] callRes;
  logic [67:0] gzdLLzicase16056;
  logic [7:0] callResR1;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLzicase16053 = {binOpR1[255:128] < binOpR1[127:0], arg1, arg2};
  zdLLzicase16053  zdLLzicase16053 (gzdLLzicase16053[66:3], gzdLLzicase16053[2:0], callRes);
  assign gzdLLzicase16056 = {binOp[255:128] < binOp[127:0], arg0, arg2};
  zdLLzicase16056  zdLLzicase16056 (gzdLLzicase16056[66:3], gzdLLzicase16056[2:0], callResR1);
  assign res = (gzdLLzicase16056[67] == 1'h1) ? callResR1 : callRes;
endmodule

module zdLLzilambda16070 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [67:0] gzdLLzicase16063;
  logic [7:0] callRes;
  logic [67:0] gzdLLzicase16066;
  logic [7:0] callResR1;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLzicase16063 = {binOpR1[255:128] < binOpR1[127:0], arg1, arg2};
  zdLLzicase16063  zdLLzicase16063 (gzdLLzicase16063[66:3], gzdLLzicase16063[2:0], callRes);
  assign gzdLLzicase16066 = {binOp[255:128] < binOp[127:0], arg0, arg2};
  zdLLzicase16066  zdLLzicase16066 (gzdLLzicase16066[66:3], gzdLLzicase16066[2:0], callResR1);
  assign res = (gzdLLzicase16066[67] == 1'h1) ? callResR1 : callRes;
endmodule

module zdLLzilambda16082 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [131:0] gzdLLzicase16074;
  logic [130:0] gzdLLzilambda16070;
  logic [7:0] callRes;
  logic [130:0] gzdLLzilambda16070R1;
  logic [7:0] callResR1;
  logic [130:0] gzdLLzilambda16070R2;
  logic [7:0] callResR2;
  logic [130:0] gzdLLzilambda16070R3;
  logic [7:0] callResR3;
  logic [130:0] gzdLLzilambda16070R4;
  logic [7:0] callResR4;
  logic [130:0] gzdLLzilambda16070R5;
  logic [7:0] callResR5;
  logic [130:0] gzdLLzilambda16070R6;
  logic [7:0] callResR6;
  logic [130:0] gzdLLzilambda16070R7;
  logic [7:0] callResR7;
  logic [63:0] resizzeR2;
  logic [2:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR6;
  logic [2:0] resizzeR7;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [127:0] resizzeR8;
  logic [131:0] gzdLLzicase16078;
  logic [130:0] gzdLLzilambda16060;
  logic [7:0] callResR8;
  logic [130:0] gzdLLzilambda16060R1;
  logic [7:0] callResR9;
  logic [130:0] gzdLLzilambda16060R2;
  logic [7:0] callResR10;
  logic [130:0] gzdLLzilambda16060R3;
  logic [7:0] callResR11;
  logic [130:0] gzdLLzilambda16060R4;
  logic [7:0] callResR12;
  logic [130:0] gzdLLzilambda16060R5;
  logic [7:0] callResR13;
  logic [130:0] gzdLLzilambda16060R6;
  logic [7:0] callResR14;
  logic [130:0] gzdLLzilambda16060R7;
  logic [7:0] callResR15;
  logic [63:0] resizzeR9;
  logic [2:0] resizzeR10;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [127:0] resizzeR11;
  logic [2:0] resizzeR12;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [255:0] binOpR14;
  logic [255:0] binOpR15;
  logic [127:0] resizzeR13;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLzicase16074 = {binOpR1[255:128] < binOpR1[127:0], arg0, arg1, arg2};
  assign gzdLLzilambda16070 = {gzdLLzicase16074[130:67], gzdLLzicase16074[66:3], 3'h0};
  zdLLzilambda16070  zdLLzilambda16070 (gzdLLzilambda16070[130:67], gzdLLzilambda16070[66:3], gzdLLzilambda16070[2:0], callRes);
  assign gzdLLzilambda16070R1 = {gzdLLzicase16074[130:67], gzdLLzicase16074[66:3], 3'h1};
  zdLLzilambda16070  zdLLzilambda16070R1 (gzdLLzilambda16070R1[130:67], gzdLLzilambda16070R1[66:3], gzdLLzilambda16070R1[2:0], callResR1);
  assign gzdLLzilambda16070R2 = {gzdLLzicase16074[130:67], gzdLLzicase16074[66:3], 3'h2};
  zdLLzilambda16070  zdLLzilambda16070R2 (gzdLLzilambda16070R2[130:67], gzdLLzilambda16070R2[66:3], gzdLLzilambda16070R2[2:0], callResR2);
  assign gzdLLzilambda16070R3 = {gzdLLzicase16074[130:67], gzdLLzicase16074[66:3], 3'h3};
  zdLLzilambda16070  zdLLzilambda16070R3 (gzdLLzilambda16070R3[130:67], gzdLLzilambda16070R3[66:3], gzdLLzilambda16070R3[2:0], callResR3);
  assign gzdLLzilambda16070R4 = {gzdLLzicase16074[130:67], gzdLLzicase16074[66:3], 3'h4};
  zdLLzilambda16070  zdLLzilambda16070R4 (gzdLLzilambda16070R4[130:67], gzdLLzilambda16070R4[66:3], gzdLLzilambda16070R4[2:0], callResR4);
  assign gzdLLzilambda16070R5 = {gzdLLzicase16074[130:67], gzdLLzicase16074[66:3], 3'h5};
  zdLLzilambda16070  zdLLzilambda16070R5 (gzdLLzilambda16070R5[130:67], gzdLLzilambda16070R5[66:3], gzdLLzilambda16070R5[2:0], callResR5);
  assign gzdLLzilambda16070R6 = {gzdLLzicase16074[130:67], gzdLLzicase16074[66:3], 3'h6};
  zdLLzilambda16070  zdLLzilambda16070R6 (gzdLLzilambda16070R6[130:67], gzdLLzilambda16070R6[66:3], gzdLLzilambda16070R6[2:0], callResR6);
  assign gzdLLzilambda16070R7 = {gzdLLzicase16074[130:67], gzdLLzicase16074[66:3], 3'h7};
  zdLLzilambda16070  zdLLzilambda16070R7 (gzdLLzilambda16070R7[130:67], gzdLLzilambda16070R7[66:3], gzdLLzilambda16070R7[2:0], callResR7);
  assign resizzeR2 = {callRes, callResR1, callResR2, callResR3, callResR4, callResR5, callResR6, callResR7};
  assign resizzeR3 = gzdLLzicase16074[2:0];
  assign binOpR2 = {128'(resizzeR3[2:0]), 128'h00000000000000000000000000000003};
  assign binOpR3 = {binOpR2[255:128] - binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[2:0];
  assign binOpR4 = {128'(resizzeR5[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR5 = {binOpR4[255:128] * binOpR4[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR6 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR7 = resizzeR6[2:0];
  assign binOpR6 = {128'h00000000000000000000000000000008, 128'(resizzeR7[2:0])};
  assign binOpR7 = {binOpR6[255:128] - binOpR6[127:0], 128'h00000000000000000000000000000001};
  assign binOpR8 = {binOpR7[255:128] - binOpR7[127:0], 128'h00000000000000000000000000000008};
  assign binOpR9 = {128'(resizzeR2[63:0]), binOpR8[255:128] * binOpR8[127:0]};
  assign resizzeR8 = binOpR9[255:128] >> binOpR9[127:0];
  assign gzdLLzicase16078 = {binOp[255:128] < binOp[127:0], arg0, arg1, arg2};
  assign gzdLLzilambda16060 = {gzdLLzicase16078[130:67], gzdLLzicase16078[66:3], 3'h0};
  zdLLzilambda16060  zdLLzilambda16060 (gzdLLzilambda16060[130:67], gzdLLzilambda16060[66:3], gzdLLzilambda16060[2:0], callResR8);
  assign gzdLLzilambda16060R1 = {gzdLLzicase16078[130:67], gzdLLzicase16078[66:3], 3'h1};
  zdLLzilambda16060  zdLLzilambda16060R1 (gzdLLzilambda16060R1[130:67], gzdLLzilambda16060R1[66:3], gzdLLzilambda16060R1[2:0], callResR9);
  assign gzdLLzilambda16060R2 = {gzdLLzicase16078[130:67], gzdLLzicase16078[66:3], 3'h2};
  zdLLzilambda16060  zdLLzilambda16060R2 (gzdLLzilambda16060R2[130:67], gzdLLzilambda16060R2[66:3], gzdLLzilambda16060R2[2:0], callResR10);
  assign gzdLLzilambda16060R3 = {gzdLLzicase16078[130:67], gzdLLzicase16078[66:3], 3'h3};
  zdLLzilambda16060  zdLLzilambda16060R3 (gzdLLzilambda16060R3[130:67], gzdLLzilambda16060R3[66:3], gzdLLzilambda16060R3[2:0], callResR11);
  assign gzdLLzilambda16060R4 = {gzdLLzicase16078[130:67], gzdLLzicase16078[66:3], 3'h4};
  zdLLzilambda16060  zdLLzilambda16060R4 (gzdLLzilambda16060R4[130:67], gzdLLzilambda16060R4[66:3], gzdLLzilambda16060R4[2:0], callResR12);
  assign gzdLLzilambda16060R5 = {gzdLLzicase16078[130:67], gzdLLzicase16078[66:3], 3'h5};
  zdLLzilambda16060  zdLLzilambda16060R5 (gzdLLzilambda16060R5[130:67], gzdLLzilambda16060R5[66:3], gzdLLzilambda16060R5[2:0], callResR13);
  assign gzdLLzilambda16060R6 = {gzdLLzicase16078[130:67], gzdLLzicase16078[66:3], 3'h6};
  zdLLzilambda16060  zdLLzilambda16060R6 (gzdLLzilambda16060R6[130:67], gzdLLzilambda16060R6[66:3], gzdLLzilambda16060R6[2:0], callResR14);
  assign gzdLLzilambda16060R7 = {gzdLLzicase16078[130:67], gzdLLzicase16078[66:3], 3'h7};
  zdLLzilambda16060  zdLLzilambda16060R7 (gzdLLzilambda16060R7[130:67], gzdLLzilambda16060R7[66:3], gzdLLzilambda16060R7[2:0], callResR15);
  assign resizzeR9 = {callResR8, callResR9, callResR10, callResR11, callResR12, callResR13, callResR14, callResR15};
  assign resizzeR10 = gzdLLzicase16078[2:0];
  assign binOpR10 = {128'(resizzeR10[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR11 = {binOpR10[255:128] * binOpR10[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR11 = binOpR11[255:128] % binOpR11[127:0];
  assign resizzeR12 = resizzeR11[2:0];
  assign binOpR12 = {128'h00000000000000000000000000000008, 128'(resizzeR12[2:0])};
  assign binOpR13 = {binOpR12[255:128] - binOpR12[127:0], 128'h00000000000000000000000000000001};
  assign binOpR14 = {binOpR13[255:128] - binOpR13[127:0], 128'h00000000000000000000000000000008};
  assign binOpR15 = {128'(resizzeR9[63:0]), binOpR14[255:128] * binOpR14[127:0]};
  assign resizzeR13 = binOpR15[255:128] >> binOpR15[127:0];
  assign res = (gzdLLzicase16078[131] == 1'h1) ? resizzeR13[7:0] : resizzeR8[7:0];
endmodule

module zdLLzilambda16092 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [67:0] gzdLLzicase16053;
  logic [7:0] callRes;
  logic [67:0] gzdLLzicase16056;
  logic [7:0] callResR1;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLzicase16053 = {binOpR1[255:128] < binOpR1[127:0], arg1, arg2};
  zdLLzicase16053  zdLLzicase16053 (gzdLLzicase16053[66:3], gzdLLzicase16053[2:0], callRes);
  assign gzdLLzicase16056 = {binOp[255:128] < binOp[127:0], arg0, arg2};
  zdLLzicase16056  zdLLzicase16056 (gzdLLzicase16056[66:3], gzdLLzicase16056[2:0], callResR1);
  assign res = (gzdLLzicase16056[67] == 1'h1) ? callResR1 : callRes;
endmodule

module zdLLzilambda16102 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [67:0] gzdLLzicase16063;
  logic [7:0] callRes;
  logic [67:0] gzdLLzicase16066;
  logic [7:0] callResR1;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLzicase16063 = {binOpR1[255:128] < binOpR1[127:0], arg1, arg2};
  zdLLzicase16063  zdLLzicase16063 (gzdLLzicase16063[66:3], gzdLLzicase16063[2:0], callRes);
  assign gzdLLzicase16066 = {binOp[255:128] < binOp[127:0], arg0, arg2};
  zdLLzicase16066  zdLLzicase16066 (gzdLLzicase16066[66:3], gzdLLzicase16066[2:0], callResR1);
  assign res = (gzdLLzicase16066[67] == 1'h1) ? callResR1 : callRes;
endmodule

module zdLLzilambda16114 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [131:0] gzdLLzicase16106;
  logic [130:0] gzdLLzilambda16102;
  logic [7:0] callRes;
  logic [130:0] gzdLLzilambda16102R1;
  logic [7:0] callResR1;
  logic [130:0] gzdLLzilambda16102R2;
  logic [7:0] callResR2;
  logic [130:0] gzdLLzilambda16102R3;
  logic [7:0] callResR3;
  logic [130:0] gzdLLzilambda16102R4;
  logic [7:0] callResR4;
  logic [130:0] gzdLLzilambda16102R5;
  logic [7:0] callResR5;
  logic [130:0] gzdLLzilambda16102R6;
  logic [7:0] callResR6;
  logic [130:0] gzdLLzilambda16102R7;
  logic [7:0] callResR7;
  logic [63:0] resizzeR2;
  logic [2:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR6;
  logic [2:0] resizzeR7;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [127:0] resizzeR8;
  logic [2:0] resizzeR9;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [127:0] resizzeR10;
  logic [131:0] gzdLLzicase16110;
  logic [130:0] gzdLLzilambda16092;
  logic [7:0] callResR8;
  logic [130:0] gzdLLzilambda16092R1;
  logic [7:0] callResR9;
  logic [130:0] gzdLLzilambda16092R2;
  logic [7:0] callResR10;
  logic [130:0] gzdLLzilambda16092R3;
  logic [7:0] callResR11;
  logic [130:0] gzdLLzilambda16092R4;
  logic [7:0] callResR12;
  logic [130:0] gzdLLzilambda16092R5;
  logic [7:0] callResR13;
  logic [130:0] gzdLLzilambda16092R6;
  logic [7:0] callResR14;
  logic [130:0] gzdLLzilambda16092R7;
  logic [7:0] callResR15;
  logic [63:0] resizzeR11;
  logic [2:0] resizzeR12;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [127:0] resizzeR13;
  logic [2:0] resizzeR14;
  logic [255:0] binOpR14;
  logic [255:0] binOpR15;
  logic [127:0] resizzeR15;
  logic [2:0] resizzeR16;
  logic [255:0] binOpR16;
  logic [255:0] binOpR17;
  logic [255:0] binOpR18;
  logic [255:0] binOpR19;
  logic [127:0] resizzeR17;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLzicase16106 = {binOpR1[255:128] < binOpR1[127:0], arg0, arg1, arg2};
  assign gzdLLzilambda16102 = {gzdLLzicase16106[130:67], gzdLLzicase16106[66:3], 3'h0};
  zdLLzilambda16102  zdLLzilambda16102 (gzdLLzilambda16102[130:67], gzdLLzilambda16102[66:3], gzdLLzilambda16102[2:0], callRes);
  assign gzdLLzilambda16102R1 = {gzdLLzicase16106[130:67], gzdLLzicase16106[66:3], 3'h1};
  zdLLzilambda16102  zdLLzilambda16102R1 (gzdLLzilambda16102R1[130:67], gzdLLzilambda16102R1[66:3], gzdLLzilambda16102R1[2:0], callResR1);
  assign gzdLLzilambda16102R2 = {gzdLLzicase16106[130:67], gzdLLzicase16106[66:3], 3'h2};
  zdLLzilambda16102  zdLLzilambda16102R2 (gzdLLzilambda16102R2[130:67], gzdLLzilambda16102R2[66:3], gzdLLzilambda16102R2[2:0], callResR2);
  assign gzdLLzilambda16102R3 = {gzdLLzicase16106[130:67], gzdLLzicase16106[66:3], 3'h3};
  zdLLzilambda16102  zdLLzilambda16102R3 (gzdLLzilambda16102R3[130:67], gzdLLzilambda16102R3[66:3], gzdLLzilambda16102R3[2:0], callResR3);
  assign gzdLLzilambda16102R4 = {gzdLLzicase16106[130:67], gzdLLzicase16106[66:3], 3'h4};
  zdLLzilambda16102  zdLLzilambda16102R4 (gzdLLzilambda16102R4[130:67], gzdLLzilambda16102R4[66:3], gzdLLzilambda16102R4[2:0], callResR4);
  assign gzdLLzilambda16102R5 = {gzdLLzicase16106[130:67], gzdLLzicase16106[66:3], 3'h5};
  zdLLzilambda16102  zdLLzilambda16102R5 (gzdLLzilambda16102R5[130:67], gzdLLzilambda16102R5[66:3], gzdLLzilambda16102R5[2:0], callResR5);
  assign gzdLLzilambda16102R6 = {gzdLLzicase16106[130:67], gzdLLzicase16106[66:3], 3'h6};
  zdLLzilambda16102  zdLLzilambda16102R6 (gzdLLzilambda16102R6[130:67], gzdLLzilambda16102R6[66:3], gzdLLzilambda16102R6[2:0], callResR6);
  assign gzdLLzilambda16102R7 = {gzdLLzicase16106[130:67], gzdLLzicase16106[66:3], 3'h7};
  zdLLzilambda16102  zdLLzilambda16102R7 (gzdLLzilambda16102R7[130:67], gzdLLzilambda16102R7[66:3], gzdLLzilambda16102R7[2:0], callResR7);
  assign resizzeR2 = {callRes, callResR1, callResR2, callResR3, callResR4, callResR5, callResR6, callResR7};
  assign resizzeR3 = gzdLLzicase16106[2:0];
  assign binOpR2 = {128'(resizzeR3[2:0]), 128'h00000000000000000000000000000003};
  assign binOpR3 = {binOpR2[255:128] - binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[2:0];
  assign binOpR4 = {128'(resizzeR5[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR5 = {binOpR4[255:128] * binOpR4[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR6 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR7 = resizzeR6[2:0];
  assign binOpR6 = {128'(resizzeR7[2:0]), 128'h00000000000000000000000000000001};
  assign binOpR7 = {binOpR6[255:128] + binOpR6[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR8 = binOpR7[255:128] % binOpR7[127:0];
  assign resizzeR9 = resizzeR8[2:0];
  assign binOpR8 = {128'h00000000000000000000000000000008, 128'(resizzeR9[2:0])};
  assign binOpR9 = {binOpR8[255:128] - binOpR8[127:0], 128'h00000000000000000000000000000001};
  assign binOpR10 = {binOpR9[255:128] - binOpR9[127:0], 128'h00000000000000000000000000000008};
  assign binOpR11 = {128'(resizzeR2[63:0]), binOpR10[255:128] * binOpR10[127:0]};
  assign resizzeR10 = binOpR11[255:128] >> binOpR11[127:0];
  assign gzdLLzicase16110 = {binOp[255:128] < binOp[127:0], arg0, arg1, arg2};
  assign gzdLLzilambda16092 = {gzdLLzicase16110[130:67], gzdLLzicase16110[66:3], 3'h0};
  zdLLzilambda16092  zdLLzilambda16092 (gzdLLzilambda16092[130:67], gzdLLzilambda16092[66:3], gzdLLzilambda16092[2:0], callResR8);
  assign gzdLLzilambda16092R1 = {gzdLLzicase16110[130:67], gzdLLzicase16110[66:3], 3'h1};
  zdLLzilambda16092  zdLLzilambda16092R1 (gzdLLzilambda16092R1[130:67], gzdLLzilambda16092R1[66:3], gzdLLzilambda16092R1[2:0], callResR9);
  assign gzdLLzilambda16092R2 = {gzdLLzicase16110[130:67], gzdLLzicase16110[66:3], 3'h2};
  zdLLzilambda16092  zdLLzilambda16092R2 (gzdLLzilambda16092R2[130:67], gzdLLzilambda16092R2[66:3], gzdLLzilambda16092R2[2:0], callResR10);
  assign gzdLLzilambda16092R3 = {gzdLLzicase16110[130:67], gzdLLzicase16110[66:3], 3'h3};
  zdLLzilambda16092  zdLLzilambda16092R3 (gzdLLzilambda16092R3[130:67], gzdLLzilambda16092R3[66:3], gzdLLzilambda16092R3[2:0], callResR11);
  assign gzdLLzilambda16092R4 = {gzdLLzicase16110[130:67], gzdLLzicase16110[66:3], 3'h4};
  zdLLzilambda16092  zdLLzilambda16092R4 (gzdLLzilambda16092R4[130:67], gzdLLzilambda16092R4[66:3], gzdLLzilambda16092R4[2:0], callResR12);
  assign gzdLLzilambda16092R5 = {gzdLLzicase16110[130:67], gzdLLzicase16110[66:3], 3'h5};
  zdLLzilambda16092  zdLLzilambda16092R5 (gzdLLzilambda16092R5[130:67], gzdLLzilambda16092R5[66:3], gzdLLzilambda16092R5[2:0], callResR13);
  assign gzdLLzilambda16092R6 = {gzdLLzicase16110[130:67], gzdLLzicase16110[66:3], 3'h6};
  zdLLzilambda16092  zdLLzilambda16092R6 (gzdLLzilambda16092R6[130:67], gzdLLzilambda16092R6[66:3], gzdLLzilambda16092R6[2:0], callResR14);
  assign gzdLLzilambda16092R7 = {gzdLLzicase16110[130:67], gzdLLzicase16110[66:3], 3'h7};
  zdLLzilambda16092  zdLLzilambda16092R7 (gzdLLzilambda16092R7[130:67], gzdLLzilambda16092R7[66:3], gzdLLzilambda16092R7[2:0], callResR15);
  assign resizzeR11 = {callResR8, callResR9, callResR10, callResR11, callResR12, callResR13, callResR14, callResR15};
  assign resizzeR12 = gzdLLzicase16110[2:0];
  assign binOpR12 = {128'(resizzeR12[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR13 = {binOpR12[255:128] * binOpR12[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR13 = binOpR13[255:128] % binOpR13[127:0];
  assign resizzeR14 = resizzeR13[2:0];
  assign binOpR14 = {128'(resizzeR14[2:0]), 128'h00000000000000000000000000000001};
  assign binOpR15 = {binOpR14[255:128] + binOpR14[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR15 = binOpR15[255:128] % binOpR15[127:0];
  assign resizzeR16 = resizzeR15[2:0];
  assign binOpR16 = {128'h00000000000000000000000000000008, 128'(resizzeR16[2:0])};
  assign binOpR17 = {binOpR16[255:128] - binOpR16[127:0], 128'h00000000000000000000000000000001};
  assign binOpR18 = {binOpR17[255:128] - binOpR17[127:0], 128'h00000000000000000000000000000008};
  assign binOpR19 = {128'(resizzeR11[63:0]), binOpR18[255:128] * binOpR18[127:0]};
  assign resizzeR17 = binOpR19[255:128] >> binOpR19[127:0];
  assign res = (gzdLLzicase16110[131] == 1'h1) ? resizzeR17[7:0] : resizzeR10[7:0];
endmodule

module zdLLzilambda16126 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [127:0] resizzeR1;
  logic [0:0] msbit;
  logic [0:0] gReWireziPreludezinot;
  logic [0:0] callRes;
  logic [2:0] resizzeR2;
  logic [127:0] resizzeR3;
  logic [0:0] msbitR1;
  logic [0:0] gReWireziPreludezinotR1;
  logic [0:0] callResR1;
  logic [131:0] gzdLLzicase16118;
  logic [130:0] gzdLLzilambda16114;
  logic [7:0] callResR2;
  logic [130:0] gzdLLzilambda16114R1;
  logic [7:0] callResR3;
  logic [130:0] gzdLLzilambda16114R2;
  logic [7:0] callResR4;
  logic [130:0] gzdLLzilambda16114R3;
  logic [7:0] callResR5;
  logic [130:0] gzdLLzilambda16114R4;
  logic [7:0] callResR6;
  logic [130:0] gzdLLzilambda16114R5;
  logic [7:0] callResR7;
  logic [130:0] gzdLLzilambda16114R6;
  logic [7:0] callResR8;
  logic [130:0] gzdLLzilambda16114R7;
  logic [7:0] callResR9;
  logic [63:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOp;
  logic [255:0] binOpR1;
  logic [127:0] resizzeR6;
  logic [2:0] resizzeR7;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR8;
  logic [2:0] resizzeR9;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [127:0] resizzeR10;
  logic [131:0] gzdLLzicase16122;
  logic [130:0] gzdLLzilambda16082;
  logic [7:0] callResR10;
  logic [130:0] gzdLLzilambda16082R1;
  logic [7:0] callResR11;
  logic [130:0] gzdLLzilambda16082R2;
  logic [7:0] callResR12;
  logic [130:0] gzdLLzilambda16082R3;
  logic [7:0] callResR13;
  logic [130:0] gzdLLzilambda16082R4;
  logic [7:0] callResR14;
  logic [130:0] gzdLLzilambda16082R5;
  logic [7:0] callResR15;
  logic [130:0] gzdLLzilambda16082R6;
  logic [7:0] callResR16;
  logic [130:0] gzdLLzilambda16082R7;
  logic [7:0] callResR17;
  logic [63:0] resizzeR11;
  logic [2:0] resizzeR12;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [127:0] resizzeR13;
  logic [2:0] resizzeR14;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [127:0] resizzeR15;
  assign resizze = arg2;
  assign resizzeR1 = 128'(resizze[2:0]);
  assign msbit = resizzeR1[0];
  assign gReWireziPreludezinot = msbit[0];
  ReWireziPreludezinot  ReWireziPreludezinot (gReWireziPreludezinot[0], callRes);
  assign resizzeR2 = arg2;
  assign resizzeR3 = 128'(resizzeR2[2:0]);
  assign msbitR1 = resizzeR3[0];
  assign gReWireziPreludezinotR1 = msbitR1[0];
  ReWireziPreludezinot  ReWireziPreludezinotR1 (gReWireziPreludezinotR1[0], callResR1);
  assign gzdLLzicase16118 = {callResR1, arg0, arg1, arg2};
  assign gzdLLzilambda16114 = {gzdLLzicase16118[130:67], gzdLLzicase16118[66:3], 3'h0};
  zdLLzilambda16114  zdLLzilambda16114 (gzdLLzilambda16114[130:67], gzdLLzilambda16114[66:3], gzdLLzilambda16114[2:0], callResR2);
  assign gzdLLzilambda16114R1 = {gzdLLzicase16118[130:67], gzdLLzicase16118[66:3], 3'h1};
  zdLLzilambda16114  zdLLzilambda16114R1 (gzdLLzilambda16114R1[130:67], gzdLLzilambda16114R1[66:3], gzdLLzilambda16114R1[2:0], callResR3);
  assign gzdLLzilambda16114R2 = {gzdLLzicase16118[130:67], gzdLLzicase16118[66:3], 3'h2};
  zdLLzilambda16114  zdLLzilambda16114R2 (gzdLLzilambda16114R2[130:67], gzdLLzilambda16114R2[66:3], gzdLLzilambda16114R2[2:0], callResR4);
  assign gzdLLzilambda16114R3 = {gzdLLzicase16118[130:67], gzdLLzicase16118[66:3], 3'h3};
  zdLLzilambda16114  zdLLzilambda16114R3 (gzdLLzilambda16114R3[130:67], gzdLLzilambda16114R3[66:3], gzdLLzilambda16114R3[2:0], callResR5);
  assign gzdLLzilambda16114R4 = {gzdLLzicase16118[130:67], gzdLLzicase16118[66:3], 3'h4};
  zdLLzilambda16114  zdLLzilambda16114R4 (gzdLLzilambda16114R4[130:67], gzdLLzilambda16114R4[66:3], gzdLLzilambda16114R4[2:0], callResR6);
  assign gzdLLzilambda16114R5 = {gzdLLzicase16118[130:67], gzdLLzicase16118[66:3], 3'h5};
  zdLLzilambda16114  zdLLzilambda16114R5 (gzdLLzilambda16114R5[130:67], gzdLLzilambda16114R5[66:3], gzdLLzilambda16114R5[2:0], callResR7);
  assign gzdLLzilambda16114R6 = {gzdLLzicase16118[130:67], gzdLLzicase16118[66:3], 3'h6};
  zdLLzilambda16114  zdLLzilambda16114R6 (gzdLLzilambda16114R6[130:67], gzdLLzilambda16114R6[66:3], gzdLLzilambda16114R6[2:0], callResR8);
  assign gzdLLzilambda16114R7 = {gzdLLzicase16118[130:67], gzdLLzicase16118[66:3], 3'h7};
  zdLLzilambda16114  zdLLzilambda16114R7 (gzdLLzilambda16114R7[130:67], gzdLLzilambda16114R7[66:3], gzdLLzilambda16114R7[2:0], callResR9);
  assign resizzeR4 = {callResR2, callResR3, callResR4, callResR5, callResR6, callResR7, callResR8, callResR9};
  assign resizzeR5 = gzdLLzicase16118[2:0];
  assign binOp = {128'(resizzeR5[2:0]), 128'h00000000000000000000000000000001};
  assign binOpR1 = {binOp[255:128] - binOp[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR6 = binOpR1[255:128] % binOpR1[127:0];
  assign resizzeR7 = resizzeR6[2:0];
  assign binOpR2 = {128'(resizzeR7[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR3 = {binOpR2[255:128] / binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR8 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR9 = resizzeR8[2:0];
  assign binOpR4 = {128'h00000000000000000000000000000008, 128'(resizzeR9[2:0])};
  assign binOpR5 = {binOpR4[255:128] - binOpR4[127:0], 128'h00000000000000000000000000000001};
  assign binOpR6 = {binOpR5[255:128] - binOpR5[127:0], 128'h00000000000000000000000000000008};
  assign binOpR7 = {128'(resizzeR4[63:0]), binOpR6[255:128] * binOpR6[127:0]};
  assign resizzeR10 = binOpR7[255:128] >> binOpR7[127:0];
  assign gzdLLzicase16122 = {callRes, arg0, arg1, arg2};
  assign gzdLLzilambda16082 = {gzdLLzicase16122[130:67], gzdLLzicase16122[66:3], 3'h0};
  zdLLzilambda16082  zdLLzilambda16082 (gzdLLzilambda16082[130:67], gzdLLzilambda16082[66:3], gzdLLzilambda16082[2:0], callResR10);
  assign gzdLLzilambda16082R1 = {gzdLLzicase16122[130:67], gzdLLzicase16122[66:3], 3'h1};
  zdLLzilambda16082  zdLLzilambda16082R1 (gzdLLzilambda16082R1[130:67], gzdLLzilambda16082R1[66:3], gzdLLzilambda16082R1[2:0], callResR11);
  assign gzdLLzilambda16082R2 = {gzdLLzicase16122[130:67], gzdLLzicase16122[66:3], 3'h2};
  zdLLzilambda16082  zdLLzilambda16082R2 (gzdLLzilambda16082R2[130:67], gzdLLzilambda16082R2[66:3], gzdLLzilambda16082R2[2:0], callResR12);
  assign gzdLLzilambda16082R3 = {gzdLLzicase16122[130:67], gzdLLzicase16122[66:3], 3'h3};
  zdLLzilambda16082  zdLLzilambda16082R3 (gzdLLzilambda16082R3[130:67], gzdLLzilambda16082R3[66:3], gzdLLzilambda16082R3[2:0], callResR13);
  assign gzdLLzilambda16082R4 = {gzdLLzicase16122[130:67], gzdLLzicase16122[66:3], 3'h4};
  zdLLzilambda16082  zdLLzilambda16082R4 (gzdLLzilambda16082R4[130:67], gzdLLzilambda16082R4[66:3], gzdLLzilambda16082R4[2:0], callResR14);
  assign gzdLLzilambda16082R5 = {gzdLLzicase16122[130:67], gzdLLzicase16122[66:3], 3'h5};
  zdLLzilambda16082  zdLLzilambda16082R5 (gzdLLzilambda16082R5[130:67], gzdLLzilambda16082R5[66:3], gzdLLzilambda16082R5[2:0], callResR15);
  assign gzdLLzilambda16082R6 = {gzdLLzicase16122[130:67], gzdLLzicase16122[66:3], 3'h6};
  zdLLzilambda16082  zdLLzilambda16082R6 (gzdLLzilambda16082R6[130:67], gzdLLzilambda16082R6[66:3], gzdLLzilambda16082R6[2:0], callResR16);
  assign gzdLLzilambda16082R7 = {gzdLLzicase16122[130:67], gzdLLzicase16122[66:3], 3'h7};
  zdLLzilambda16082  zdLLzilambda16082R7 (gzdLLzilambda16082R7[130:67], gzdLLzilambda16082R7[66:3], gzdLLzilambda16082R7[2:0], callResR17);
  assign resizzeR11 = {callResR10, callResR11, callResR12, callResR13, callResR14, callResR15, callResR16, callResR17};
  assign resizzeR12 = gzdLLzicase16122[2:0];
  assign binOpR8 = {128'(resizzeR12[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR9 = {binOpR8[255:128] / binOpR8[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR13 = binOpR9[255:128] % binOpR9[127:0];
  assign resizzeR14 = resizzeR13[2:0];
  assign binOpR10 = {128'h00000000000000000000000000000008, 128'(resizzeR14[2:0])};
  assign binOpR11 = {binOpR10[255:128] - binOpR10[127:0], 128'h00000000000000000000000000000001};
  assign binOpR12 = {binOpR11[255:128] - binOpR11[127:0], 128'h00000000000000000000000000000008};
  assign binOpR13 = {128'(resizzeR11[63:0]), binOpR12[255:128] * binOpR12[127:0]};
  assign resizzeR15 = binOpR13[255:128] >> binOpR13[127:0];
  assign res = (gzdLLzicase16122[131] == 1'h1) ? resizzeR15[7:0] : resizzeR10[7:0];
endmodule

module zdLLzilambda16136 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [67:0] gzdLLzicase16053;
  logic [7:0] callRes;
  logic [67:0] gzdLLzicase16056;
  logic [7:0] callResR1;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLzicase16053 = {binOpR1[255:128] < binOpR1[127:0], arg1, arg2};
  zdLLzicase16053  zdLLzicase16053 (gzdLLzicase16053[66:3], gzdLLzicase16053[2:0], callRes);
  assign gzdLLzicase16056 = {binOp[255:128] < binOp[127:0], arg0, arg2};
  zdLLzicase16056  zdLLzicase16056 (gzdLLzicase16056[66:3], gzdLLzicase16056[2:0], callResR1);
  assign res = (gzdLLzicase16056[67] == 1'h1) ? callResR1 : callRes;
endmodule

module zdLLzilambda16146 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [67:0] gzdLLzicase16063;
  logic [7:0] callRes;
  logic [67:0] gzdLLzicase16066;
  logic [7:0] callResR1;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLzicase16063 = {binOpR1[255:128] < binOpR1[127:0], arg1, arg2};
  zdLLzicase16063  zdLLzicase16063 (gzdLLzicase16063[66:3], gzdLLzicase16063[2:0], callRes);
  assign gzdLLzicase16066 = {binOp[255:128] < binOp[127:0], arg0, arg2};
  zdLLzicase16066  zdLLzicase16066 (gzdLLzicase16066[66:3], gzdLLzicase16066[2:0], callResR1);
  assign res = (gzdLLzicase16066[67] == 1'h1) ? callResR1 : callRes;
endmodule

module zdLLzilambda16158 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [131:0] gzdLLzicase16150;
  logic [130:0] gzdLLzilambda16146;
  logic [7:0] callRes;
  logic [130:0] gzdLLzilambda16146R1;
  logic [7:0] callResR1;
  logic [130:0] gzdLLzilambda16146R2;
  logic [7:0] callResR2;
  logic [130:0] gzdLLzilambda16146R3;
  logic [7:0] callResR3;
  logic [130:0] gzdLLzilambda16146R4;
  logic [7:0] callResR4;
  logic [130:0] gzdLLzilambda16146R5;
  logic [7:0] callResR5;
  logic [130:0] gzdLLzilambda16146R6;
  logic [7:0] callResR6;
  logic [130:0] gzdLLzilambda16146R7;
  logic [7:0] callResR7;
  logic [63:0] resizzeR2;
  logic [2:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR6;
  logic [2:0] resizzeR7;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [127:0] resizzeR8;
  logic [131:0] gzdLLzicase16154;
  logic [130:0] gzdLLzilambda16136;
  logic [7:0] callResR8;
  logic [130:0] gzdLLzilambda16136R1;
  logic [7:0] callResR9;
  logic [130:0] gzdLLzilambda16136R2;
  logic [7:0] callResR10;
  logic [130:0] gzdLLzilambda16136R3;
  logic [7:0] callResR11;
  logic [130:0] gzdLLzilambda16136R4;
  logic [7:0] callResR12;
  logic [130:0] gzdLLzilambda16136R5;
  logic [7:0] callResR13;
  logic [130:0] gzdLLzilambda16136R6;
  logic [7:0] callResR14;
  logic [130:0] gzdLLzilambda16136R7;
  logic [7:0] callResR15;
  logic [63:0] resizzeR9;
  logic [2:0] resizzeR10;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [127:0] resizzeR11;
  logic [2:0] resizzeR12;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [255:0] binOpR14;
  logic [255:0] binOpR15;
  logic [127:0] resizzeR13;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLzicase16150 = {binOpR1[255:128] < binOpR1[127:0], arg0, arg1, arg2};
  assign gzdLLzilambda16146 = {gzdLLzicase16150[130:67], gzdLLzicase16150[66:3], 3'h0};
  zdLLzilambda16146  zdLLzilambda16146 (gzdLLzilambda16146[130:67], gzdLLzilambda16146[66:3], gzdLLzilambda16146[2:0], callRes);
  assign gzdLLzilambda16146R1 = {gzdLLzicase16150[130:67], gzdLLzicase16150[66:3], 3'h1};
  zdLLzilambda16146  zdLLzilambda16146R1 (gzdLLzilambda16146R1[130:67], gzdLLzilambda16146R1[66:3], gzdLLzilambda16146R1[2:0], callResR1);
  assign gzdLLzilambda16146R2 = {gzdLLzicase16150[130:67], gzdLLzicase16150[66:3], 3'h2};
  zdLLzilambda16146  zdLLzilambda16146R2 (gzdLLzilambda16146R2[130:67], gzdLLzilambda16146R2[66:3], gzdLLzilambda16146R2[2:0], callResR2);
  assign gzdLLzilambda16146R3 = {gzdLLzicase16150[130:67], gzdLLzicase16150[66:3], 3'h3};
  zdLLzilambda16146  zdLLzilambda16146R3 (gzdLLzilambda16146R3[130:67], gzdLLzilambda16146R3[66:3], gzdLLzilambda16146R3[2:0], callResR3);
  assign gzdLLzilambda16146R4 = {gzdLLzicase16150[130:67], gzdLLzicase16150[66:3], 3'h4};
  zdLLzilambda16146  zdLLzilambda16146R4 (gzdLLzilambda16146R4[130:67], gzdLLzilambda16146R4[66:3], gzdLLzilambda16146R4[2:0], callResR4);
  assign gzdLLzilambda16146R5 = {gzdLLzicase16150[130:67], gzdLLzicase16150[66:3], 3'h5};
  zdLLzilambda16146  zdLLzilambda16146R5 (gzdLLzilambda16146R5[130:67], gzdLLzilambda16146R5[66:3], gzdLLzilambda16146R5[2:0], callResR5);
  assign gzdLLzilambda16146R6 = {gzdLLzicase16150[130:67], gzdLLzicase16150[66:3], 3'h6};
  zdLLzilambda16146  zdLLzilambda16146R6 (gzdLLzilambda16146R6[130:67], gzdLLzilambda16146R6[66:3], gzdLLzilambda16146R6[2:0], callResR6);
  assign gzdLLzilambda16146R7 = {gzdLLzicase16150[130:67], gzdLLzicase16150[66:3], 3'h7};
  zdLLzilambda16146  zdLLzilambda16146R7 (gzdLLzilambda16146R7[130:67], gzdLLzilambda16146R7[66:3], gzdLLzilambda16146R7[2:0], callResR7);
  assign resizzeR2 = {callRes, callResR1, callResR2, callResR3, callResR4, callResR5, callResR6, callResR7};
  assign resizzeR3 = gzdLLzicase16150[2:0];
  assign binOpR2 = {128'(resizzeR3[2:0]), 128'h00000000000000000000000000000003};
  assign binOpR3 = {binOpR2[255:128] - binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[2:0];
  assign binOpR4 = {128'(resizzeR5[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR5 = {binOpR4[255:128] * binOpR4[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR6 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR7 = resizzeR6[2:0];
  assign binOpR6 = {128'h00000000000000000000000000000008, 128'(resizzeR7[2:0])};
  assign binOpR7 = {binOpR6[255:128] - binOpR6[127:0], 128'h00000000000000000000000000000001};
  assign binOpR8 = {binOpR7[255:128] - binOpR7[127:0], 128'h00000000000000000000000000000008};
  assign binOpR9 = {128'(resizzeR2[63:0]), binOpR8[255:128] * binOpR8[127:0]};
  assign resizzeR8 = binOpR9[255:128] >> binOpR9[127:0];
  assign gzdLLzicase16154 = {binOp[255:128] < binOp[127:0], arg0, arg1, arg2};
  assign gzdLLzilambda16136 = {gzdLLzicase16154[130:67], gzdLLzicase16154[66:3], 3'h0};
  zdLLzilambda16136  zdLLzilambda16136 (gzdLLzilambda16136[130:67], gzdLLzilambda16136[66:3], gzdLLzilambda16136[2:0], callResR8);
  assign gzdLLzilambda16136R1 = {gzdLLzicase16154[130:67], gzdLLzicase16154[66:3], 3'h1};
  zdLLzilambda16136  zdLLzilambda16136R1 (gzdLLzilambda16136R1[130:67], gzdLLzilambda16136R1[66:3], gzdLLzilambda16136R1[2:0], callResR9);
  assign gzdLLzilambda16136R2 = {gzdLLzicase16154[130:67], gzdLLzicase16154[66:3], 3'h2};
  zdLLzilambda16136  zdLLzilambda16136R2 (gzdLLzilambda16136R2[130:67], gzdLLzilambda16136R2[66:3], gzdLLzilambda16136R2[2:0], callResR10);
  assign gzdLLzilambda16136R3 = {gzdLLzicase16154[130:67], gzdLLzicase16154[66:3], 3'h3};
  zdLLzilambda16136  zdLLzilambda16136R3 (gzdLLzilambda16136R3[130:67], gzdLLzilambda16136R3[66:3], gzdLLzilambda16136R3[2:0], callResR11);
  assign gzdLLzilambda16136R4 = {gzdLLzicase16154[130:67], gzdLLzicase16154[66:3], 3'h4};
  zdLLzilambda16136  zdLLzilambda16136R4 (gzdLLzilambda16136R4[130:67], gzdLLzilambda16136R4[66:3], gzdLLzilambda16136R4[2:0], callResR12);
  assign gzdLLzilambda16136R5 = {gzdLLzicase16154[130:67], gzdLLzicase16154[66:3], 3'h5};
  zdLLzilambda16136  zdLLzilambda16136R5 (gzdLLzilambda16136R5[130:67], gzdLLzilambda16136R5[66:3], gzdLLzilambda16136R5[2:0], callResR13);
  assign gzdLLzilambda16136R6 = {gzdLLzicase16154[130:67], gzdLLzicase16154[66:3], 3'h6};
  zdLLzilambda16136  zdLLzilambda16136R6 (gzdLLzilambda16136R6[130:67], gzdLLzilambda16136R6[66:3], gzdLLzilambda16136R6[2:0], callResR14);
  assign gzdLLzilambda16136R7 = {gzdLLzicase16154[130:67], gzdLLzicase16154[66:3], 3'h7};
  zdLLzilambda16136  zdLLzilambda16136R7 (gzdLLzilambda16136R7[130:67], gzdLLzilambda16136R7[66:3], gzdLLzilambda16136R7[2:0], callResR15);
  assign resizzeR9 = {callResR8, callResR9, callResR10, callResR11, callResR12, callResR13, callResR14, callResR15};
  assign resizzeR10 = gzdLLzicase16154[2:0];
  assign binOpR10 = {128'(resizzeR10[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR11 = {binOpR10[255:128] * binOpR10[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR11 = binOpR11[255:128] % binOpR11[127:0];
  assign resizzeR12 = resizzeR11[2:0];
  assign binOpR12 = {128'h00000000000000000000000000000008, 128'(resizzeR12[2:0])};
  assign binOpR13 = {binOpR12[255:128] - binOpR12[127:0], 128'h00000000000000000000000000000001};
  assign binOpR14 = {binOpR13[255:128] - binOpR13[127:0], 128'h00000000000000000000000000000008};
  assign binOpR15 = {128'(resizzeR9[63:0]), binOpR14[255:128] * binOpR14[127:0]};
  assign resizzeR13 = binOpR15[255:128] >> binOpR15[127:0];
  assign res = (gzdLLzicase16154[131] == 1'h1) ? resizzeR13[7:0] : resizzeR8[7:0];
endmodule

module zdLLzilambda16168 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [67:0] gzdLLzicase16053;
  logic [7:0] callRes;
  logic [67:0] gzdLLzicase16056;
  logic [7:0] callResR1;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLzicase16053 = {binOpR1[255:128] < binOpR1[127:0], arg1, arg2};
  zdLLzicase16053  zdLLzicase16053 (gzdLLzicase16053[66:3], gzdLLzicase16053[2:0], callRes);
  assign gzdLLzicase16056 = {binOp[255:128] < binOp[127:0], arg0, arg2};
  zdLLzicase16056  zdLLzicase16056 (gzdLLzicase16056[66:3], gzdLLzicase16056[2:0], callResR1);
  assign res = (gzdLLzicase16056[67] == 1'h1) ? callResR1 : callRes;
endmodule

module zdLLzilambda16178 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [67:0] gzdLLzicase16063;
  logic [7:0] callRes;
  logic [67:0] gzdLLzicase16066;
  logic [7:0] callResR1;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLzicase16063 = {binOpR1[255:128] < binOpR1[127:0], arg1, arg2};
  zdLLzicase16063  zdLLzicase16063 (gzdLLzicase16063[66:3], gzdLLzicase16063[2:0], callRes);
  assign gzdLLzicase16066 = {binOp[255:128] < binOp[127:0], arg0, arg2};
  zdLLzicase16066  zdLLzicase16066 (gzdLLzicase16066[66:3], gzdLLzicase16066[2:0], callResR1);
  assign res = (gzdLLzicase16066[67] == 1'h1) ? callResR1 : callRes;
endmodule

module zdLLzilambda16190 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [131:0] gzdLLzicase16182;
  logic [130:0] gzdLLzilambda16178;
  logic [7:0] callRes;
  logic [130:0] gzdLLzilambda16178R1;
  logic [7:0] callResR1;
  logic [130:0] gzdLLzilambda16178R2;
  logic [7:0] callResR2;
  logic [130:0] gzdLLzilambda16178R3;
  logic [7:0] callResR3;
  logic [130:0] gzdLLzilambda16178R4;
  logic [7:0] callResR4;
  logic [130:0] gzdLLzilambda16178R5;
  logic [7:0] callResR5;
  logic [130:0] gzdLLzilambda16178R6;
  logic [7:0] callResR6;
  logic [130:0] gzdLLzilambda16178R7;
  logic [7:0] callResR7;
  logic [63:0] resizzeR2;
  logic [2:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR6;
  logic [2:0] resizzeR7;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [127:0] resizzeR8;
  logic [2:0] resizzeR9;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [127:0] resizzeR10;
  logic [131:0] gzdLLzicase16186;
  logic [130:0] gzdLLzilambda16168;
  logic [7:0] callResR8;
  logic [130:0] gzdLLzilambda16168R1;
  logic [7:0] callResR9;
  logic [130:0] gzdLLzilambda16168R2;
  logic [7:0] callResR10;
  logic [130:0] gzdLLzilambda16168R3;
  logic [7:0] callResR11;
  logic [130:0] gzdLLzilambda16168R4;
  logic [7:0] callResR12;
  logic [130:0] gzdLLzilambda16168R5;
  logic [7:0] callResR13;
  logic [130:0] gzdLLzilambda16168R6;
  logic [7:0] callResR14;
  logic [130:0] gzdLLzilambda16168R7;
  logic [7:0] callResR15;
  logic [63:0] resizzeR11;
  logic [2:0] resizzeR12;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [127:0] resizzeR13;
  logic [2:0] resizzeR14;
  logic [255:0] binOpR14;
  logic [255:0] binOpR15;
  logic [127:0] resizzeR15;
  logic [2:0] resizzeR16;
  logic [255:0] binOpR16;
  logic [255:0] binOpR17;
  logic [255:0] binOpR18;
  logic [255:0] binOpR19;
  logic [127:0] resizzeR17;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLzicase16182 = {binOpR1[255:128] < binOpR1[127:0], arg0, arg1, arg2};
  assign gzdLLzilambda16178 = {gzdLLzicase16182[130:67], gzdLLzicase16182[66:3], 3'h0};
  zdLLzilambda16178  zdLLzilambda16178 (gzdLLzilambda16178[130:67], gzdLLzilambda16178[66:3], gzdLLzilambda16178[2:0], callRes);
  assign gzdLLzilambda16178R1 = {gzdLLzicase16182[130:67], gzdLLzicase16182[66:3], 3'h1};
  zdLLzilambda16178  zdLLzilambda16178R1 (gzdLLzilambda16178R1[130:67], gzdLLzilambda16178R1[66:3], gzdLLzilambda16178R1[2:0], callResR1);
  assign gzdLLzilambda16178R2 = {gzdLLzicase16182[130:67], gzdLLzicase16182[66:3], 3'h2};
  zdLLzilambda16178  zdLLzilambda16178R2 (gzdLLzilambda16178R2[130:67], gzdLLzilambda16178R2[66:3], gzdLLzilambda16178R2[2:0], callResR2);
  assign gzdLLzilambda16178R3 = {gzdLLzicase16182[130:67], gzdLLzicase16182[66:3], 3'h3};
  zdLLzilambda16178  zdLLzilambda16178R3 (gzdLLzilambda16178R3[130:67], gzdLLzilambda16178R3[66:3], gzdLLzilambda16178R3[2:0], callResR3);
  assign gzdLLzilambda16178R4 = {gzdLLzicase16182[130:67], gzdLLzicase16182[66:3], 3'h4};
  zdLLzilambda16178  zdLLzilambda16178R4 (gzdLLzilambda16178R4[130:67], gzdLLzilambda16178R4[66:3], gzdLLzilambda16178R4[2:0], callResR4);
  assign gzdLLzilambda16178R5 = {gzdLLzicase16182[130:67], gzdLLzicase16182[66:3], 3'h5};
  zdLLzilambda16178  zdLLzilambda16178R5 (gzdLLzilambda16178R5[130:67], gzdLLzilambda16178R5[66:3], gzdLLzilambda16178R5[2:0], callResR5);
  assign gzdLLzilambda16178R6 = {gzdLLzicase16182[130:67], gzdLLzicase16182[66:3], 3'h6};
  zdLLzilambda16178  zdLLzilambda16178R6 (gzdLLzilambda16178R6[130:67], gzdLLzilambda16178R6[66:3], gzdLLzilambda16178R6[2:0], callResR6);
  assign gzdLLzilambda16178R7 = {gzdLLzicase16182[130:67], gzdLLzicase16182[66:3], 3'h7};
  zdLLzilambda16178  zdLLzilambda16178R7 (gzdLLzilambda16178R7[130:67], gzdLLzilambda16178R7[66:3], gzdLLzilambda16178R7[2:0], callResR7);
  assign resizzeR2 = {callRes, callResR1, callResR2, callResR3, callResR4, callResR5, callResR6, callResR7};
  assign resizzeR3 = gzdLLzicase16182[2:0];
  assign binOpR2 = {128'(resizzeR3[2:0]), 128'h00000000000000000000000000000003};
  assign binOpR3 = {binOpR2[255:128] - binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[2:0];
  assign binOpR4 = {128'(resizzeR5[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR5 = {binOpR4[255:128] * binOpR4[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR6 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR7 = resizzeR6[2:0];
  assign binOpR6 = {128'(resizzeR7[2:0]), 128'h00000000000000000000000000000001};
  assign binOpR7 = {binOpR6[255:128] + binOpR6[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR8 = binOpR7[255:128] % binOpR7[127:0];
  assign resizzeR9 = resizzeR8[2:0];
  assign binOpR8 = {128'h00000000000000000000000000000008, 128'(resizzeR9[2:0])};
  assign binOpR9 = {binOpR8[255:128] - binOpR8[127:0], 128'h00000000000000000000000000000001};
  assign binOpR10 = {binOpR9[255:128] - binOpR9[127:0], 128'h00000000000000000000000000000008};
  assign binOpR11 = {128'(resizzeR2[63:0]), binOpR10[255:128] * binOpR10[127:0]};
  assign resizzeR10 = binOpR11[255:128] >> binOpR11[127:0];
  assign gzdLLzicase16186 = {binOp[255:128] < binOp[127:0], arg0, arg1, arg2};
  assign gzdLLzilambda16168 = {gzdLLzicase16186[130:67], gzdLLzicase16186[66:3], 3'h0};
  zdLLzilambda16168  zdLLzilambda16168 (gzdLLzilambda16168[130:67], gzdLLzilambda16168[66:3], gzdLLzilambda16168[2:0], callResR8);
  assign gzdLLzilambda16168R1 = {gzdLLzicase16186[130:67], gzdLLzicase16186[66:3], 3'h1};
  zdLLzilambda16168  zdLLzilambda16168R1 (gzdLLzilambda16168R1[130:67], gzdLLzilambda16168R1[66:3], gzdLLzilambda16168R1[2:0], callResR9);
  assign gzdLLzilambda16168R2 = {gzdLLzicase16186[130:67], gzdLLzicase16186[66:3], 3'h2};
  zdLLzilambda16168  zdLLzilambda16168R2 (gzdLLzilambda16168R2[130:67], gzdLLzilambda16168R2[66:3], gzdLLzilambda16168R2[2:0], callResR10);
  assign gzdLLzilambda16168R3 = {gzdLLzicase16186[130:67], gzdLLzicase16186[66:3], 3'h3};
  zdLLzilambda16168  zdLLzilambda16168R3 (gzdLLzilambda16168R3[130:67], gzdLLzilambda16168R3[66:3], gzdLLzilambda16168R3[2:0], callResR11);
  assign gzdLLzilambda16168R4 = {gzdLLzicase16186[130:67], gzdLLzicase16186[66:3], 3'h4};
  zdLLzilambda16168  zdLLzilambda16168R4 (gzdLLzilambda16168R4[130:67], gzdLLzilambda16168R4[66:3], gzdLLzilambda16168R4[2:0], callResR12);
  assign gzdLLzilambda16168R5 = {gzdLLzicase16186[130:67], gzdLLzicase16186[66:3], 3'h5};
  zdLLzilambda16168  zdLLzilambda16168R5 (gzdLLzilambda16168R5[130:67], gzdLLzilambda16168R5[66:3], gzdLLzilambda16168R5[2:0], callResR13);
  assign gzdLLzilambda16168R6 = {gzdLLzicase16186[130:67], gzdLLzicase16186[66:3], 3'h6};
  zdLLzilambda16168  zdLLzilambda16168R6 (gzdLLzilambda16168R6[130:67], gzdLLzilambda16168R6[66:3], gzdLLzilambda16168R6[2:0], callResR14);
  assign gzdLLzilambda16168R7 = {gzdLLzicase16186[130:67], gzdLLzicase16186[66:3], 3'h7};
  zdLLzilambda16168  zdLLzilambda16168R7 (gzdLLzilambda16168R7[130:67], gzdLLzilambda16168R7[66:3], gzdLLzilambda16168R7[2:0], callResR15);
  assign resizzeR11 = {callResR8, callResR9, callResR10, callResR11, callResR12, callResR13, callResR14, callResR15};
  assign resizzeR12 = gzdLLzicase16186[2:0];
  assign binOpR12 = {128'(resizzeR12[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR13 = {binOpR12[255:128] * binOpR12[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR13 = binOpR13[255:128] % binOpR13[127:0];
  assign resizzeR14 = resizzeR13[2:0];
  assign binOpR14 = {128'(resizzeR14[2:0]), 128'h00000000000000000000000000000001};
  assign binOpR15 = {binOpR14[255:128] + binOpR14[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR15 = binOpR15[255:128] % binOpR15[127:0];
  assign resizzeR16 = resizzeR15[2:0];
  assign binOpR16 = {128'h00000000000000000000000000000008, 128'(resizzeR16[2:0])};
  assign binOpR17 = {binOpR16[255:128] - binOpR16[127:0], 128'h00000000000000000000000000000001};
  assign binOpR18 = {binOpR17[255:128] - binOpR17[127:0], 128'h00000000000000000000000000000008};
  assign binOpR19 = {128'(resizzeR11[63:0]), binOpR18[255:128] * binOpR18[127:0]};
  assign resizzeR17 = binOpR19[255:128] >> binOpR19[127:0];
  assign res = (gzdLLzicase16186[131] == 1'h1) ? resizzeR17[7:0] : resizzeR10[7:0];
endmodule

module zdLLzilambda16202 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [127:0] resizzeR1;
  logic [0:0] msbit;
  logic [0:0] gReWireziPreludezinot;
  logic [0:0] callRes;
  logic [2:0] resizzeR2;
  logic [127:0] resizzeR3;
  logic [0:0] msbitR1;
  logic [0:0] gReWireziPreludezinotR1;
  logic [0:0] callResR1;
  logic [131:0] gzdLLzicase16194;
  logic [130:0] gzdLLzilambda16190;
  logic [7:0] callResR2;
  logic [130:0] gzdLLzilambda16190R1;
  logic [7:0] callResR3;
  logic [130:0] gzdLLzilambda16190R2;
  logic [7:0] callResR4;
  logic [130:0] gzdLLzilambda16190R3;
  logic [7:0] callResR5;
  logic [130:0] gzdLLzilambda16190R4;
  logic [7:0] callResR6;
  logic [130:0] gzdLLzilambda16190R5;
  logic [7:0] callResR7;
  logic [130:0] gzdLLzilambda16190R6;
  logic [7:0] callResR8;
  logic [130:0] gzdLLzilambda16190R7;
  logic [7:0] callResR9;
  logic [63:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOp;
  logic [255:0] binOpR1;
  logic [127:0] resizzeR6;
  logic [2:0] resizzeR7;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR8;
  logic [2:0] resizzeR9;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR10;
  logic [2:0] resizzeR11;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [127:0] resizzeR12;
  logic [131:0] gzdLLzicase16198;
  logic [130:0] gzdLLzilambda16158;
  logic [7:0] callResR10;
  logic [130:0] gzdLLzilambda16158R1;
  logic [7:0] callResR11;
  logic [130:0] gzdLLzilambda16158R2;
  logic [7:0] callResR12;
  logic [130:0] gzdLLzilambda16158R3;
  logic [7:0] callResR13;
  logic [130:0] gzdLLzilambda16158R4;
  logic [7:0] callResR14;
  logic [130:0] gzdLLzilambda16158R5;
  logic [7:0] callResR15;
  logic [130:0] gzdLLzilambda16158R6;
  logic [7:0] callResR16;
  logic [130:0] gzdLLzilambda16158R7;
  logic [7:0] callResR17;
  logic [63:0] resizzeR13;
  logic [2:0] resizzeR14;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [127:0] resizzeR15;
  logic [2:0] resizzeR16;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [127:0] resizzeR17;
  logic [2:0] resizzeR18;
  logic [255:0] binOpR14;
  logic [255:0] binOpR15;
  logic [255:0] binOpR16;
  logic [255:0] binOpR17;
  logic [127:0] resizzeR19;
  assign resizze = arg2;
  assign resizzeR1 = 128'(resizze[2:0]);
  assign msbit = resizzeR1[0];
  assign gReWireziPreludezinot = msbit[0];
  ReWireziPreludezinot  ReWireziPreludezinot (gReWireziPreludezinot[0], callRes);
  assign resizzeR2 = arg2;
  assign resizzeR3 = 128'(resizzeR2[2:0]);
  assign msbitR1 = resizzeR3[0];
  assign gReWireziPreludezinotR1 = msbitR1[0];
  ReWireziPreludezinot  ReWireziPreludezinotR1 (gReWireziPreludezinotR1[0], callResR1);
  assign gzdLLzicase16194 = {callResR1, arg0, arg1, arg2};
  assign gzdLLzilambda16190 = {gzdLLzicase16194[130:67], gzdLLzicase16194[66:3], 3'h0};
  zdLLzilambda16190  zdLLzilambda16190 (gzdLLzilambda16190[130:67], gzdLLzilambda16190[66:3], gzdLLzilambda16190[2:0], callResR2);
  assign gzdLLzilambda16190R1 = {gzdLLzicase16194[130:67], gzdLLzicase16194[66:3], 3'h1};
  zdLLzilambda16190  zdLLzilambda16190R1 (gzdLLzilambda16190R1[130:67], gzdLLzilambda16190R1[66:3], gzdLLzilambda16190R1[2:0], callResR3);
  assign gzdLLzilambda16190R2 = {gzdLLzicase16194[130:67], gzdLLzicase16194[66:3], 3'h2};
  zdLLzilambda16190  zdLLzilambda16190R2 (gzdLLzilambda16190R2[130:67], gzdLLzilambda16190R2[66:3], gzdLLzilambda16190R2[2:0], callResR4);
  assign gzdLLzilambda16190R3 = {gzdLLzicase16194[130:67], gzdLLzicase16194[66:3], 3'h3};
  zdLLzilambda16190  zdLLzilambda16190R3 (gzdLLzilambda16190R3[130:67], gzdLLzilambda16190R3[66:3], gzdLLzilambda16190R3[2:0], callResR5);
  assign gzdLLzilambda16190R4 = {gzdLLzicase16194[130:67], gzdLLzicase16194[66:3], 3'h4};
  zdLLzilambda16190  zdLLzilambda16190R4 (gzdLLzilambda16190R4[130:67], gzdLLzilambda16190R4[66:3], gzdLLzilambda16190R4[2:0], callResR6);
  assign gzdLLzilambda16190R5 = {gzdLLzicase16194[130:67], gzdLLzicase16194[66:3], 3'h5};
  zdLLzilambda16190  zdLLzilambda16190R5 (gzdLLzilambda16190R5[130:67], gzdLLzilambda16190R5[66:3], gzdLLzilambda16190R5[2:0], callResR7);
  assign gzdLLzilambda16190R6 = {gzdLLzicase16194[130:67], gzdLLzicase16194[66:3], 3'h6};
  zdLLzilambda16190  zdLLzilambda16190R6 (gzdLLzilambda16190R6[130:67], gzdLLzilambda16190R6[66:3], gzdLLzilambda16190R6[2:0], callResR8);
  assign gzdLLzilambda16190R7 = {gzdLLzicase16194[130:67], gzdLLzicase16194[66:3], 3'h7};
  zdLLzilambda16190  zdLLzilambda16190R7 (gzdLLzilambda16190R7[130:67], gzdLLzilambda16190R7[66:3], gzdLLzilambda16190R7[2:0], callResR9);
  assign resizzeR4 = {callResR2, callResR3, callResR4, callResR5, callResR6, callResR7, callResR8, callResR9};
  assign resizzeR5 = gzdLLzicase16194[2:0];
  assign binOp = {128'(resizzeR5[2:0]), 128'h00000000000000000000000000000001};
  assign binOpR1 = {binOp[255:128] - binOp[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR6 = binOpR1[255:128] % binOpR1[127:0];
  assign resizzeR7 = resizzeR6[2:0];
  assign binOpR2 = {128'h00000000000000000000000000000003, 128'(resizzeR7[2:0])};
  assign binOpR3 = {binOpR2[255:128] + binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR8 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR9 = resizzeR8[2:0];
  assign binOpR4 = {128'(resizzeR9[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR5 = {binOpR4[255:128] / binOpR4[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR10 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR11 = resizzeR10[2:0];
  assign binOpR6 = {128'h00000000000000000000000000000008, 128'(resizzeR11[2:0])};
  assign binOpR7 = {binOpR6[255:128] - binOpR6[127:0], 128'h00000000000000000000000000000001};
  assign binOpR8 = {binOpR7[255:128] - binOpR7[127:0], 128'h00000000000000000000000000000008};
  assign binOpR9 = {128'(resizzeR4[63:0]), binOpR8[255:128] * binOpR8[127:0]};
  assign resizzeR12 = binOpR9[255:128] >> binOpR9[127:0];
  assign gzdLLzicase16198 = {callRes, arg0, arg1, arg2};
  assign gzdLLzilambda16158 = {gzdLLzicase16198[130:67], gzdLLzicase16198[66:3], 3'h0};
  zdLLzilambda16158  zdLLzilambda16158 (gzdLLzilambda16158[130:67], gzdLLzilambda16158[66:3], gzdLLzilambda16158[2:0], callResR10);
  assign gzdLLzilambda16158R1 = {gzdLLzicase16198[130:67], gzdLLzicase16198[66:3], 3'h1};
  zdLLzilambda16158  zdLLzilambda16158R1 (gzdLLzilambda16158R1[130:67], gzdLLzilambda16158R1[66:3], gzdLLzilambda16158R1[2:0], callResR11);
  assign gzdLLzilambda16158R2 = {gzdLLzicase16198[130:67], gzdLLzicase16198[66:3], 3'h2};
  zdLLzilambda16158  zdLLzilambda16158R2 (gzdLLzilambda16158R2[130:67], gzdLLzilambda16158R2[66:3], gzdLLzilambda16158R2[2:0], callResR12);
  assign gzdLLzilambda16158R3 = {gzdLLzicase16198[130:67], gzdLLzicase16198[66:3], 3'h3};
  zdLLzilambda16158  zdLLzilambda16158R3 (gzdLLzilambda16158R3[130:67], gzdLLzilambda16158R3[66:3], gzdLLzilambda16158R3[2:0], callResR13);
  assign gzdLLzilambda16158R4 = {gzdLLzicase16198[130:67], gzdLLzicase16198[66:3], 3'h4};
  zdLLzilambda16158  zdLLzilambda16158R4 (gzdLLzilambda16158R4[130:67], gzdLLzilambda16158R4[66:3], gzdLLzilambda16158R4[2:0], callResR14);
  assign gzdLLzilambda16158R5 = {gzdLLzicase16198[130:67], gzdLLzicase16198[66:3], 3'h5};
  zdLLzilambda16158  zdLLzilambda16158R5 (gzdLLzilambda16158R5[130:67], gzdLLzilambda16158R5[66:3], gzdLLzilambda16158R5[2:0], callResR15);
  assign gzdLLzilambda16158R6 = {gzdLLzicase16198[130:67], gzdLLzicase16198[66:3], 3'h6};
  zdLLzilambda16158  zdLLzilambda16158R6 (gzdLLzilambda16158R6[130:67], gzdLLzilambda16158R6[66:3], gzdLLzilambda16158R6[2:0], callResR16);
  assign gzdLLzilambda16158R7 = {gzdLLzicase16198[130:67], gzdLLzicase16198[66:3], 3'h7};
  zdLLzilambda16158  zdLLzilambda16158R7 (gzdLLzilambda16158R7[130:67], gzdLLzilambda16158R7[66:3], gzdLLzilambda16158R7[2:0], callResR17);
  assign resizzeR13 = {callResR10, callResR11, callResR12, callResR13, callResR14, callResR15, callResR16, callResR17};
  assign resizzeR14 = gzdLLzicase16198[2:0];
  assign binOpR10 = {128'h00000000000000000000000000000003, 128'(resizzeR14[2:0])};
  assign binOpR11 = {binOpR10[255:128] + binOpR10[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR15 = binOpR11[255:128] % binOpR11[127:0];
  assign resizzeR16 = resizzeR15[2:0];
  assign binOpR12 = {128'(resizzeR16[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR13 = {binOpR12[255:128] / binOpR12[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR17 = binOpR13[255:128] % binOpR13[127:0];
  assign resizzeR18 = resizzeR17[2:0];
  assign binOpR14 = {128'h00000000000000000000000000000008, 128'(resizzeR18[2:0])};
  assign binOpR15 = {binOpR14[255:128] - binOpR14[127:0], 128'h00000000000000000000000000000001};
  assign binOpR16 = {binOpR15[255:128] - binOpR15[127:0], 128'h00000000000000000000000000000008};
  assign binOpR17 = {128'(resizzeR13[63:0]), binOpR16[255:128] * binOpR16[127:0]};
  assign resizzeR19 = binOpR17[255:128] >> binOpR17[127:0];
  assign res = (gzdLLzicase16198[131] == 1'h1) ? resizzeR19[7:0] : resizzeR12[7:0];
endmodule

module ReWireziPreludezinot (input logic [0:0] arg0,
  output logic [0:0] res);
  logic [0:0] lit;
  assign lit = arg0;
  assign res = (lit[0] == 1'h1) ? 1'h0 : 1'h1;
endmodule