module test1 (input logic [31:0] a, input logic [31:0] b, output logic out);
      assign out = a[0] & b[0];
endmodule

module test2 (input logic [31:0] a, input logic [31:0] b, output logic out);
      assign out = a[0] & b[0];
endmodule

module test3 (input logic [31:0] a, input logic [31:0] b, output logic out);
      assign out = a[0] & b[0];
endmodule

module test4 (input logic [31:0] a, input logic [31:0] b, output logic out);
      assign out = a[0] & b[0];
endmodule

