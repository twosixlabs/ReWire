module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [0:0] __in0,
  input logic [31:0] __in1,
  output logic [0:0] __out0,
  output logic [0:0] __out1);
  logic [71:0] main_repl1_in;
  logic [104:0] zll_main_repl58_in;
  logic [71:0] zll_main_repl15_in;
  logic [71:0] zll_main_repl94_in;
  logic [80:0] zll_main_repl94_out;
  logic [71:0] zll_main_repl113_in;
  logic [70:0] zll_main_repl30_in;
  logic [70:0] zll_main_repl74_in;
  logic [77:0] zll_main_repl11_in;
  logic [77:0] zll_main_repl68_in;
  logic [112:0] zll_main_repl47_in;
  logic [112:0] zll_main_repl109_in;
  logic [109:0] zll_main_repl96_in;
  logic [109:0] zll_main_repl79_in;
  logic [109:0] zll_main_repl42_in;
  logic [109:0] zll_main_repl102_in;
  logic [109:0] zll_main_repl3_in;
  logic [77:0] zll_main_repl103_in;
  logic [84:0] zll_main_repl82_in;
  logic [84:0] zll_main_repl99_in;
  logic [84:0] zll_main_repl52_in;
  logic [84:0] zll_main_repl23_in;
  logic [84:0] zll_main_repl95_in;
  logic [84:0] zll_main_repl112_in;
  logic [77:0] zll_main_repl14_in;
  logic [38:0] main_nextpc_in;
  logic [38:0] main_nextpc_out;
  logic [38:0] zll_main_repl110_in;
  logic [80:0] zll_main_repl110_out;
  logic [80:0] zll_main_repl101_in;
  logic [80:0] zll_main_repl101_out;
  logic [77:0] zll_main_repl57_in;
  logic [70:0] zll_main_repl93_in;
  logic [70:0] zll_main_repl107_in;
  logic [38:0] main_getreg_in;
  logic [70:0] main_getreg_out;
  logic [70:0] zll_main_repl85_in;
  logic [80:0] zll_main_repl85_out;
  logic [112:0] zll_main_repl40_in;
  logic [112:0] zll_main_repl51_in;
  logic [102:0] zll_main_repl61_in;
  logic [63:0] test4_in;
  logic [0:0] extres;
  logic [77:0] zll_main_repl83_in;
  logic [70:0] zll_main_repl18_in;
  logic [70:0] zll_main_repl88_in;
  logic [38:0] main_getreg_inR1;
  logic [70:0] main_getreg_outR1;
  logic [70:0] zll_main_repl85_inR1;
  logic [80:0] zll_main_repl85_outR1;
  logic [112:0] zll_main_repl111_in;
  logic [112:0] zll_main_repl38_in;
  logic [102:0] zll_main_repl100_in;
  logic [63:0] test3_in;
  logic [0:0] extresR1;
  logic [77:0] zll_main_repl87_in;
  logic [70:0] zll_main_repl62_in;
  logic [70:0] zll_main_repl36_in;
  logic [38:0] main_getreg_inR2;
  logic [70:0] main_getreg_outR2;
  logic [70:0] zll_main_repl85_inR2;
  logic [80:0] zll_main_repl85_outR2;
  logic [112:0] zll_main_repl60_in;
  logic [112:0] zll_main_repl86_in;
  logic [102:0] zll_main_repl108_in;
  logic [63:0] test2_in;
  logic [0:0] extresR2;
  logic [77:0] zll_main_repl98_in;
  logic [80:0] zll_main_repl98_out;
  logic [77:0] zll_main_repl48_in;
  logic [80:0] zll_main_repl48_out;
  logic [77:0] zll_main_repl98_inR1;
  logic [80:0] zll_main_repl98_outR1;
  logic [77:0] zll_main_repl48_inR1;
  logic [80:0] zll_main_repl48_outR1;
  logic [39:0] __padding;
  logic [31:0] __st0;
  logic [6:0] __st1;
  logic [31:0] __st0_next;
  logic [6:0] __st1_next;
  assign main_repl1_in = {{__in0, __in1}, {__st0, __st1}};
  assign zll_main_repl58_in = {main_repl1_in[71:39], main_repl1_in[71:39], main_repl1_in[38:0]};
  assign zll_main_repl15_in = {zll_main_repl58_in[104:72], zll_main_repl58_in[38:0]};
  assign zll_main_repl94_in = {zll_main_repl15_in[38:0], zll_main_repl15_in[71:39]};
  ZLL_Main_repl94  inst (zll_main_repl94_in[71:33], zll_main_repl94_out);
  assign zll_main_repl113_in = {zll_main_repl58_in[38:0], zll_main_repl58_in[71:39]};
  assign zll_main_repl30_in = {zll_main_repl113_in[71:33], zll_main_repl113_in[31:0]};
  assign zll_main_repl74_in = {zll_main_repl30_in[31:0], zll_main_repl30_in[70:32]};
  assign zll_main_repl11_in = {zll_main_repl74_in[38:0], zll_main_repl74_in[38:0]};
  assign zll_main_repl68_in = zll_main_repl11_in[77:0];
  assign zll_main_repl47_in = {zll_main_repl74_in[70:39], {3'h2, zll_main_repl68_in[77:39], zll_main_repl68_in[38:0]}};
  assign zll_main_repl109_in = {zll_main_repl47_in[112:81], zll_main_repl47_in[80:0]};
  assign zll_main_repl96_in = {zll_main_repl109_in[112:81], zll_main_repl109_in[77:39], zll_main_repl109_in[38:0]};
  assign zll_main_repl79_in = {zll_main_repl96_in[38:0], zll_main_repl96_in[109:78], zll_main_repl96_in[77:39]};
  assign zll_main_repl42_in = {zll_main_repl79_in[70:39], zll_main_repl79_in[109:71], zll_main_repl79_in[38:7], zll_main_repl79_in[6:0]};
  assign zll_main_repl102_in = {zll_main_repl42_in[109:78], zll_main_repl42_in[38:7], zll_main_repl42_in[77:39], zll_main_repl42_in[6:0]};
  assign zll_main_repl3_in = {zll_main_repl102_in[109:78], zll_main_repl102_in[77:46], zll_main_repl102_in[6:0], zll_main_repl102_in[45:7]};
  assign zll_main_repl103_in = {zll_main_repl3_in[109:78], zll_main_repl3_in[45:39], zll_main_repl3_in[38:0]};
  assign zll_main_repl82_in = {zll_main_repl103_in[77:46], zll_main_repl103_in[45:39], zll_main_repl103_in[45:39], zll_main_repl103_in[38:0]};
  assign zll_main_repl99_in = {zll_main_repl82_in[84:53], zll_main_repl82_in[52:46], zll_main_repl82_in[52:46], zll_main_repl82_in[38:0]};
  assign zll_main_repl52_in = {zll_main_repl99_in[84:53], zll_main_repl99_in[52:46], zll_main_repl99_in[52:46], zll_main_repl99_in[38:0]};
  assign zll_main_repl23_in = {zll_main_repl52_in[84:53], zll_main_repl52_in[52:46], zll_main_repl52_in[52:46], zll_main_repl52_in[38:0]};
  assign zll_main_repl95_in = {zll_main_repl23_in[84:53], zll_main_repl23_in[52:46], zll_main_repl23_in[52:46], zll_main_repl23_in[38:0]};
  assign zll_main_repl112_in = {zll_main_repl95_in[84:53], zll_main_repl95_in[52:46], zll_main_repl95_in[52:46], zll_main_repl95_in[38:0]};
  assign zll_main_repl14_in = {zll_main_repl112_in[84:53], zll_main_repl112_in[52:46], zll_main_repl112_in[38:0]};
  assign main_nextpc_in = zll_main_repl14_in[38:0];
  Main_nextPC  instR1 (main_nextpc_in[38:0], main_nextpc_out);
  assign zll_main_repl110_in = main_nextpc_out;
  ZLL_Main_repl110  instR2 (zll_main_repl110_in[38:0], zll_main_repl110_out);
  assign zll_main_repl101_in = zll_main_repl110_out;
  ZLL_Main_repl101  instR3 (zll_main_repl101_in[80:0], zll_main_repl101_out);
  assign zll_main_repl57_in = {zll_main_repl14_in[38:0], zll_main_repl14_in[77:46], zll_main_repl14_in[45:39]};
  assign zll_main_repl93_in = {zll_main_repl57_in[77:39], zll_main_repl57_in[38:7]};
  assign zll_main_repl107_in = {zll_main_repl93_in[31:0], zll_main_repl93_in[70:32]};
  assign main_getreg_in = zll_main_repl107_in[38:0];
  Main_getReg  instR4 (main_getreg_in[38:0], main_getreg_out);
  assign zll_main_repl85_in = main_getreg_out;
  ZLL_Main_repl85  instR5 (zll_main_repl85_in[70:0], zll_main_repl85_out);
  assign zll_main_repl40_in = {zll_main_repl107_in[70:39], zll_main_repl85_out};
  assign zll_main_repl51_in = {zll_main_repl40_in[112:81], zll_main_repl40_in[80:0]};
  assign zll_main_repl61_in = {zll_main_repl51_in[112:81], zll_main_repl51_in[70:39], zll_main_repl51_in[38:0]};
  assign test4_in = {zll_main_repl61_in[102:71], zll_main_repl61_in[70:39]};
  test4  instR6 (test4_in[63:32], test4_in[31:0], extres[0]);
  assign zll_main_repl83_in = {zll_main_repl112_in[38:0], zll_main_repl112_in[84:53], zll_main_repl112_in[45:39]};
  assign zll_main_repl18_in = {zll_main_repl83_in[77:39], zll_main_repl83_in[38:7]};
  assign zll_main_repl88_in = {zll_main_repl18_in[31:0], zll_main_repl18_in[70:32]};
  assign main_getreg_inR1 = zll_main_repl88_in[38:0];
  Main_getReg  instR7 (main_getreg_inR1[38:0], main_getreg_outR1);
  assign zll_main_repl85_inR1 = main_getreg_outR1;
  ZLL_Main_repl85  instR8 (zll_main_repl85_inR1[70:0], zll_main_repl85_outR1);
  assign zll_main_repl111_in = {zll_main_repl88_in[70:39], zll_main_repl85_outR1};
  assign zll_main_repl38_in = {zll_main_repl111_in[112:81], zll_main_repl111_in[80:0]};
  assign zll_main_repl100_in = {zll_main_repl38_in[112:81], zll_main_repl38_in[70:39], zll_main_repl38_in[38:0]};
  assign test3_in = {zll_main_repl100_in[102:71], zll_main_repl100_in[70:39]};
  test3  instR9 (test3_in[63:32], test3_in[31:0], extresR1[0]);
  assign zll_main_repl87_in = {zll_main_repl95_in[38:0], zll_main_repl95_in[84:53], zll_main_repl95_in[45:39]};
  assign zll_main_repl62_in = {zll_main_repl87_in[77:39], zll_main_repl87_in[38:7]};
  assign zll_main_repl36_in = {zll_main_repl62_in[31:0], zll_main_repl62_in[70:32]};
  assign main_getreg_inR2 = zll_main_repl36_in[38:0];
  Main_getReg  instR10 (main_getreg_inR2[38:0], main_getreg_outR2);
  assign zll_main_repl85_inR2 = main_getreg_outR2;
  ZLL_Main_repl85  instR11 (zll_main_repl85_inR2[70:0], zll_main_repl85_outR2);
  assign zll_main_repl60_in = {zll_main_repl36_in[70:39], zll_main_repl85_outR2};
  assign zll_main_repl86_in = {zll_main_repl60_in[112:81], zll_main_repl60_in[80:0]};
  assign zll_main_repl108_in = {zll_main_repl86_in[112:81], zll_main_repl86_in[70:39], zll_main_repl86_in[38:0]};
  assign test2_in = {zll_main_repl108_in[102:71], zll_main_repl108_in[70:39]};
  test2  instR12 (test2_in[63:32], test2_in[31:0], extresR2[0]);
  assign zll_main_repl98_in = {zll_main_repl23_in[38:0], zll_main_repl23_in[84:53], zll_main_repl23_in[45:39]};
  ZLL_Main_repl98  instR13 (zll_main_repl98_in[77:39], zll_main_repl98_in[38:7], zll_main_repl98_out);
  assign zll_main_repl48_in = {zll_main_repl52_in[38:0], zll_main_repl52_in[84:53], zll_main_repl52_in[45:39]};
  ZLL_Main_repl48  instR14 (zll_main_repl48_in[77:39], zll_main_repl48_in[38:7], zll_main_repl48_out);
  assign zll_main_repl98_inR1 = {zll_main_repl99_in[38:0], zll_main_repl99_in[84:53], zll_main_repl99_in[45:39]};
  ZLL_Main_repl98  instR15 (zll_main_repl98_inR1[77:39], zll_main_repl98_inR1[38:7], zll_main_repl98_outR1);
  assign zll_main_repl48_inR1 = {zll_main_repl82_in[38:0], zll_main_repl82_in[84:53], zll_main_repl82_in[45:39]};
  ZLL_Main_repl48  instR16 (zll_main_repl48_inR1[77:39], zll_main_repl48_inR1[38:7], zll_main_repl48_outR1);
  assign {__padding, __out0, __out1, __st0_next, __st1_next} = (zll_main_repl113_in[32] == 1'h0) ? ((zll_main_repl48_inR1[6:0] == 7'h0) ? zll_main_repl48_outR1 : ((zll_main_repl98_inR1[6:0] == 7'h1) ? zll_main_repl98_outR1 : ((zll_main_repl48_in[6:0] == 7'h2) ? zll_main_repl48_out : ((zll_main_repl98_in[6:0] == 7'h3) ? zll_main_repl98_out : ((zll_main_repl87_in[6:0] == 7'h4) ? {{1'h1, {6'h28{1'h0}}}, extresR2, zll_main_repl108_in[38:0]} : ((zll_main_repl83_in[6:0] == 7'h5) ? {{1'h1, {6'h28{1'h0}}}, extresR1, zll_main_repl100_in[38:0]} : ((zll_main_repl57_in[6:0] == 7'h6) ? {{1'h1, {6'h28{1'h0}}}, extres, zll_main_repl61_in[38:0]} : zll_main_repl101_out))))))) : zll_main_repl94_out;
  initial {__st0, __st1} = {6'h27{1'h0}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      {__st0, __st1} <= {6'h27{1'h0}};
    end else begin
      {__st0, __st1} <= {__st0_next, __st1_next};
    end
  end
endmodule

module ZLL_Main_repl110 (input logic [38:0] arg0,
  output logic [80:0] res);
  assign res = {{3'h1, {6'h27{1'h0}}}, arg0};
endmodule

module ZLL_Main_repl101 (input logic [80:0] arg0,
  output logic [80:0] res);
  logic [80:0] zll_main_repl94_in;
  logic [80:0] zll_main_repl94_out;
  assign zll_main_repl94_in = arg0;
  ZLL_Main_repl94  inst (zll_main_repl94_in[38:0], zll_main_repl94_out);
  assign res = zll_main_repl94_out;
endmodule

module ZLL_Main_repl98 (input logic [38:0] arg0,
  input logic [31:0] arg1,
  output logic [80:0] res);
  logic [70:0] zll_main_repl105_in;
  logic [70:0] zll_main_repl65_in;
  logic [38:0] main_getreg_in;
  logic [70:0] main_getreg_out;
  logic [70:0] zll_main_repl85_in;
  logic [80:0] zll_main_repl85_out;
  logic [112:0] zll_main_repl89_in;
  logic [112:0] zll_main_repl97_in;
  logic [102:0] zll_main_repl64_in;
  logic [63:0] test1_in;
  logic [0:0] extres;
  assign zll_main_repl105_in = {arg0, arg1};
  assign zll_main_repl65_in = {zll_main_repl105_in[31:0], zll_main_repl105_in[70:32]};
  assign main_getreg_in = zll_main_repl65_in[38:0];
  Main_getReg  inst (main_getreg_in[38:0], main_getreg_out);
  assign zll_main_repl85_in = main_getreg_out;
  ZLL_Main_repl85  instR1 (zll_main_repl85_in[70:0], zll_main_repl85_out);
  assign zll_main_repl89_in = {zll_main_repl65_in[70:39], zll_main_repl85_out};
  assign zll_main_repl97_in = {zll_main_repl89_in[112:81], zll_main_repl89_in[80:0]};
  assign zll_main_repl64_in = {zll_main_repl97_in[112:81], zll_main_repl97_in[70:39], zll_main_repl97_in[38:0]};
  assign test1_in = {zll_main_repl64_in[102:71], zll_main_repl64_in[70:39]};
  test1  instR2 (test1_in[63:32], test1_in[31:0], extres[0]);
  assign res = {{1'h1, {6'h28{1'h0}}}, extres, zll_main_repl64_in[38:0]};
endmodule

module ZLL_Main_repl94 (input logic [38:0] arg0,
  output logic [80:0] res);
  logic [38:0] zll_main_repl106_in;
  assign zll_main_repl106_in = arg0;
  assign res = {42'h20000000002, zll_main_repl106_in[38:0]};
endmodule

module Main_getReg (input logic [38:0] arg0,
  output logic [70:0] res);
  logic [77:0] zll_main_getreg1_in;
  logic [77:0] zll_main_getreg3_in;
  logic [77:0] zll_main_getreg4_in;
  logic [77:0] zll_main_getreg5_in;
  logic [77:0] zll_main_getreg2_in;
  assign zll_main_getreg1_in = {arg0, arg0};
  assign zll_main_getreg3_in = zll_main_getreg1_in[77:0];
  assign zll_main_getreg4_in = {zll_main_getreg3_in[38:0], zll_main_getreg3_in[77:39]};
  assign zll_main_getreg5_in = {zll_main_getreg4_in[38:7], zll_main_getreg4_in[77:39], zll_main_getreg4_in[6:0]};
  assign zll_main_getreg2_in = {zll_main_getreg5_in[77:46], zll_main_getreg5_in[6:0], zll_main_getreg5_in[45:7]};
  assign res = {zll_main_getreg2_in[77:46], zll_main_getreg2_in[38:0]};
endmodule

module ZLL_Main_repl85 (input logic [70:0] arg0,
  output logic [80:0] res);
  logic [70:0] zll_main_repl67_in;
  assign zll_main_repl67_in = arg0;
  assign res = {10'h0, zll_main_repl67_in[70:39], zll_main_repl67_in[38:0]};
endmodule

module ZLL_Main_repl48 (input logic [38:0] arg0,
  input logic [31:0] arg1,
  output logic [80:0] res);
  logic [70:0] zll_main_repl114_in;
  logic [70:0] zll_main_repl59_in;
  logic [70:0] zll_main_putreg4_in;
  logic [109:0] zll_main_putreg9_in;
  logic [109:0] zll_main_putreg13_in;
  logic [109:0] zll_main_putreg5_in;
  logic [109:0] zll_main_putreg11_in;
  logic [109:0] zll_main_putreg3_in;
  logic [77:0] zll_main_putreg8_in;
  logic [38:0] zll_main_repl110_in;
  logic [80:0] zll_main_repl110_out;
  logic [80:0] zll_main_repl55_in;
  logic [80:0] zll_main_repl39_in;
  logic [38:0] zll_main_repl63_in;
  logic [38:0] main_nextpc_in;
  logic [38:0] main_nextpc_out;
  logic [38:0] zll_main_repl110_inR1;
  logic [80:0] zll_main_repl110_outR1;
  logic [80:0] zll_main_repl101_in;
  logic [80:0] zll_main_repl101_out;
  assign zll_main_repl114_in = {arg0, arg1};
  assign zll_main_repl59_in = {zll_main_repl114_in[31:0], zll_main_repl114_in[70:32]};
  assign zll_main_putreg4_in = {zll_main_repl59_in[70:39], zll_main_repl59_in[38:0]};
  assign zll_main_putreg9_in = {zll_main_putreg4_in[70:39], zll_main_putreg4_in[38:0], zll_main_putreg4_in[38:0]};
  assign zll_main_putreg13_in = {zll_main_putreg9_in[109:78], zll_main_putreg9_in[77:0]};
  assign zll_main_putreg5_in = {zll_main_putreg13_in[38:0], zll_main_putreg13_in[109:78], zll_main_putreg13_in[77:39]};
  assign zll_main_putreg11_in = {zll_main_putreg5_in[109:71], zll_main_putreg5_in[38:7], zll_main_putreg5_in[70:39], zll_main_putreg5_in[6:0]};
  assign zll_main_putreg3_in = {zll_main_putreg11_in[38:7], zll_main_putreg11_in[70:39], zll_main_putreg11_in[6:0], zll_main_putreg11_in[109:71]};
  assign zll_main_putreg8_in = {zll_main_putreg3_in[109:78], zll_main_putreg3_in[45:39], zll_main_putreg3_in[38:0]};
  assign zll_main_repl110_in = {zll_main_putreg8_in[77:46], zll_main_putreg8_in[45:39]};
  ZLL_Main_repl110  inst (zll_main_repl110_in[38:0], zll_main_repl110_out);
  assign zll_main_repl55_in = zll_main_repl110_out;
  assign zll_main_repl39_in = zll_main_repl55_in[80:0];
  assign zll_main_repl63_in = zll_main_repl39_in[38:0];
  assign main_nextpc_in = zll_main_repl63_in[38:0];
  Main_nextPC  instR1 (main_nextpc_in[38:0], main_nextpc_out);
  assign zll_main_repl110_inR1 = main_nextpc_out;
  ZLL_Main_repl110  instR2 (zll_main_repl110_inR1[38:0], zll_main_repl110_outR1);
  assign zll_main_repl101_in = zll_main_repl110_outR1;
  ZLL_Main_repl101  instR3 (zll_main_repl101_in[80:0], zll_main_repl101_out);
  assign res = zll_main_repl101_out;
endmodule

module Main_nextPC (input logic [38:0] arg0,
  output logic [38:0] res);
  logic [77:0] zll_main_nextpc7_in;
  logic [77:0] zll_main_nextpc5_in;
  logic [77:0] zll_main_nextpc1_in;
  logic [77:0] zll_main_nextpc3_in;
  logic [77:0] zll_main_nextpc4_in;
  logic [6:0] od19_programcounter_incpc_in;
  logic [13:0] zll_od19_programcounter_incpc213_in;
  logic [13:0] zll_od19_programcounter_incpc129_in;
  logic [13:0] zll_od19_programcounter_incpc70_in;
  logic [13:0] zll_od19_programcounter_incpc105_in;
  logic [13:0] zll_od19_programcounter_incpc2_in;
  logic [13:0] zll_od19_programcounter_incpc118_in;
  logic [13:0] zll_od19_programcounter_incpc208_in;
  logic [13:0] zll_od19_programcounter_incpc172_in;
  logic [13:0] zll_od19_programcounter_incpc98_in;
  logic [13:0] zll_od19_programcounter_incpc34_in;
  logic [13:0] zll_od19_programcounter_incpc116_in;
  logic [13:0] zll_od19_programcounter_incpc72_in;
  logic [13:0] zll_od19_programcounter_incpc4_in;
  logic [13:0] zll_od19_programcounter_incpc148_in;
  logic [13:0] zll_od19_programcounter_incpc121_in;
  logic [13:0] zll_od19_programcounter_incpc77_in;
  logic [13:0] zll_od19_programcounter_incpc12_in;
  logic [13:0] zll_od19_programcounter_incpc39_in;
  logic [13:0] zll_od19_programcounter_incpc161_in;
  logic [13:0] zll_od19_programcounter_incpc26_in;
  logic [13:0] zll_od19_programcounter_incpc111_in;
  logic [13:0] zll_od19_programcounter_incpc219_in;
  logic [13:0] zll_od19_programcounter_incpc8_in;
  logic [13:0] zll_od19_programcounter_incpc147_in;
  logic [13:0] zll_od19_programcounter_incpc60_in;
  logic [13:0] zll_od19_programcounter_incpc202_in;
  logic [13:0] zll_od19_programcounter_incpc120_in;
  logic [13:0] zll_od19_programcounter_incpc182_in;
  logic [13:0] zll_od19_programcounter_incpc114_in;
  logic [13:0] zll_od19_programcounter_incpc196_in;
  logic [13:0] zll_od19_programcounter_incpc236_in;
  logic [13:0] zll_od19_programcounter_incpc164_in;
  logic [13:0] zll_od19_programcounter_incpc226_in;
  logic [13:0] zll_od19_programcounter_incpc123_in;
  logic [13:0] zll_od19_programcounter_incpc55_in;
  logic [13:0] zll_od19_programcounter_incpc175_in;
  logic [13:0] zll_od19_programcounter_incpc224_in;
  logic [13:0] zll_od19_programcounter_incpc71_in;
  logic [13:0] zll_od19_programcounter_incpc198_in;
  logic [13:0] zll_od19_programcounter_incpc50_in;
  logic [13:0] zll_od19_programcounter_incpc128_in;
  logic [13:0] zll_od19_programcounter_incpc27_in;
  logic [13:0] zll_od19_programcounter_incpc38_in;
  logic [13:0] zll_od19_programcounter_incpc173_in;
  logic [13:0] zll_od19_programcounter_incpc117_in;
  logic [13:0] zll_od19_programcounter_incpc134_in;
  logic [13:0] zll_od19_programcounter_incpc59_in;
  logic [13:0] zll_od19_programcounter_incpc227_in;
  logic [13:0] zll_od19_programcounter_incpc183_in;
  logic [13:0] zll_od19_programcounter_incpc253_in;
  logic [13:0] zll_od19_programcounter_incpc203_in;
  logic [13:0] zll_od19_programcounter_incpc125_in;
  logic [13:0] zll_od19_programcounter_incpc144_in;
  logic [13:0] zll_od19_programcounter_incpc113_in;
  logic [13:0] zll_od19_programcounter_incpc23_in;
  logic [13:0] zll_od19_programcounter_incpc231_in;
  logic [13:0] zll_od19_programcounter_incpc212_in;
  logic [13:0] zll_od19_programcounter_incpc190_in;
  logic [13:0] zll_od19_programcounter_incpc245_in;
  logic [13:0] zll_od19_programcounter_incpc52_in;
  logic [13:0] zll_od19_programcounter_incpc56_in;
  logic [13:0] zll_od19_programcounter_incpc131_in;
  logic [13:0] zll_od19_programcounter_incpc51_in;
  logic [13:0] zll_od19_programcounter_incpc230_in;
  logic [13:0] zll_od19_programcounter_incpc168_in;
  logic [13:0] zll_od19_programcounter_incpc127_in;
  logic [13:0] zll_od19_programcounter_incpc41_in;
  logic [13:0] zll_od19_programcounter_incpc18_in;
  logic [13:0] zll_od19_programcounter_incpc174_in;
  logic [13:0] zll_od19_programcounter_incpc112_in;
  logic [13:0] zll_od19_programcounter_incpc24_in;
  logic [13:0] zll_od19_programcounter_incpc66_in;
  logic [13:0] zll_od19_programcounter_incpc35_in;
  logic [13:0] zll_od19_programcounter_incpc215_in;
  logic [13:0] zll_od19_programcounter_incpc69_in;
  logic [13:0] zll_od19_programcounter_incpc136_in;
  logic [13:0] zll_od19_programcounter_incpc187_in;
  logic [13:0] zll_od19_programcounter_incpc241_in;
  logic [13:0] zll_od19_programcounter_incpc81_in;
  logic [13:0] zll_od19_programcounter_incpc169_in;
  logic [13:0] zll_od19_programcounter_incpc207_in;
  logic [13:0] zll_od19_programcounter_incpc193_in;
  logic [13:0] zll_od19_programcounter_incpc218_in;
  logic [13:0] zll_od19_programcounter_incpc109_in;
  logic [13:0] zll_od19_programcounter_incpc156_in;
  logic [13:0] zll_od19_programcounter_incpc115_in;
  logic [13:0] zll_od19_programcounter_incpc53_in;
  logic [13:0] zll_od19_programcounter_incpc151_in;
  logic [13:0] zll_od19_programcounter_incpc63_in;
  logic [13:0] zll_od19_programcounter_incpc106_in;
  logic [13:0] zll_od19_programcounter_incpc142_in;
  logic [13:0] zll_od19_programcounter_incpc191_in;
  logic [13:0] zll_od19_programcounter_incpc204_in;
  logic [13:0] zll_od19_programcounter_incpc119_in;
  logic [13:0] zll_od19_programcounter_incpc90_in;
  logic [13:0] zll_od19_programcounter_incpc85_in;
  logic [13:0] zll_od19_programcounter_incpc62_in;
  logic [13:0] zll_od19_programcounter_incpc94_in;
  logic [13:0] zll_od19_programcounter_incpc186_in;
  logic [13:0] zll_od19_programcounter_incpc11_in;
  logic [13:0] zll_od19_programcounter_incpc37_in;
  logic [13:0] zll_od19_programcounter_incpc167_in;
  logic [13:0] zll_od19_programcounter_incpc247_in;
  logic [13:0] zll_od19_programcounter_incpc185_in;
  logic [13:0] zll_od19_programcounter_incpc80_in;
  logic [13:0] zll_od19_programcounter_incpc145_in;
  logic [13:0] zll_od19_programcounter_incpc10_in;
  logic [13:0] zll_od19_programcounter_incpc49_in;
  logic [13:0] zll_od19_programcounter_incpc93_in;
  logic [13:0] zll_od19_programcounter_incpc91_in;
  logic [13:0] zll_od19_programcounter_incpc163_in;
  logic [13:0] zll_od19_programcounter_incpc64_in;
  logic [13:0] zll_od19_programcounter_incpc101_in;
  logic [13:0] zll_od19_programcounter_incpc238_in;
  logic [13:0] zll_od19_programcounter_incpc221_in;
  logic [13:0] zll_od19_programcounter_incpc78_in;
  logic [13:0] zll_od19_programcounter_incpc22_in;
  logic [13:0] zll_od19_programcounter_incpc220_in;
  logic [13:0] zll_od19_programcounter_incpc97_in;
  logic [13:0] zll_od19_programcounter_incpc143_in;
  logic [13:0] zll_od19_programcounter_incpc197_in;
  logic [13:0] zll_od19_programcounter_incpc194_in;
  logic [13:0] zll_od19_programcounter_incpc158_in;
  logic [13:0] zll_od19_programcounter_incpc40_in;
  logic [13:0] zll_od19_programcounter_incpc250_in;
  logic [13:0] zll_od19_programcounter_incpc171_in;
  logic [6:0] lit_in;
  logic [6:0] lit_inR1;
  logic [6:0] lit_inR2;
  logic [6:0] lit_inR3;
  logic [6:0] lit_inR4;
  logic [6:0] lit_inR5;
  logic [6:0] lit_inR6;
  logic [6:0] lit_inR7;
  logic [6:0] lit_inR8;
  logic [6:0] lit_inR9;
  logic [6:0] lit_inR10;
  logic [6:0] lit_inR11;
  logic [6:0] lit_inR12;
  logic [6:0] lit_inR13;
  logic [6:0] lit_inR14;
  logic [6:0] lit_inR15;
  logic [6:0] lit_inR16;
  logic [6:0] lit_inR17;
  logic [6:0] lit_inR18;
  logic [6:0] lit_inR19;
  logic [6:0] lit_inR20;
  logic [6:0] lit_inR21;
  logic [6:0] lit_inR22;
  logic [6:0] lit_inR23;
  logic [6:0] lit_inR24;
  logic [6:0] lit_inR25;
  logic [6:0] lit_inR26;
  logic [6:0] lit_inR27;
  logic [6:0] lit_inR28;
  logic [6:0] lit_inR29;
  logic [6:0] lit_inR30;
  logic [6:0] lit_inR31;
  logic [6:0] lit_inR32;
  logic [6:0] lit_inR33;
  logic [6:0] lit_inR34;
  logic [6:0] lit_inR35;
  logic [6:0] lit_inR36;
  logic [6:0] lit_inR37;
  logic [6:0] lit_inR38;
  logic [6:0] lit_inR39;
  logic [6:0] lit_inR40;
  logic [6:0] lit_inR41;
  logic [6:0] lit_inR42;
  logic [6:0] lit_inR43;
  logic [6:0] lit_inR44;
  logic [6:0] lit_inR45;
  logic [6:0] lit_inR46;
  logic [6:0] lit_inR47;
  logic [6:0] lit_inR48;
  logic [6:0] lit_inR49;
  logic [6:0] lit_inR50;
  logic [6:0] lit_inR51;
  logic [6:0] lit_inR52;
  logic [6:0] lit_inR53;
  logic [6:0] lit_inR54;
  logic [6:0] lit_inR55;
  logic [6:0] lit_inR56;
  logic [6:0] lit_inR57;
  logic [6:0] lit_inR58;
  logic [6:0] lit_inR59;
  logic [6:0] lit_inR60;
  logic [6:0] lit_inR61;
  logic [6:0] lit_inR62;
  logic [6:0] lit_inR63;
  logic [6:0] lit_inR64;
  logic [6:0] lit_inR65;
  logic [6:0] lit_inR66;
  logic [6:0] lit_inR67;
  logic [6:0] lit_inR68;
  logic [6:0] lit_inR69;
  logic [6:0] lit_inR70;
  logic [6:0] lit_inR71;
  logic [6:0] lit_inR72;
  logic [6:0] lit_inR73;
  logic [6:0] lit_inR74;
  logic [6:0] lit_inR75;
  logic [6:0] lit_inR76;
  logic [6:0] lit_inR77;
  logic [6:0] lit_inR78;
  logic [6:0] lit_inR79;
  logic [6:0] lit_inR80;
  logic [6:0] lit_inR81;
  logic [6:0] lit_inR82;
  logic [6:0] lit_inR83;
  logic [6:0] lit_inR84;
  logic [6:0] lit_inR85;
  logic [6:0] lit_inR86;
  logic [6:0] lit_inR87;
  logic [6:0] lit_inR88;
  logic [6:0] lit_inR89;
  logic [6:0] lit_inR90;
  logic [6:0] lit_inR91;
  logic [6:0] lit_inR92;
  logic [6:0] lit_inR93;
  logic [6:0] lit_inR94;
  logic [6:0] lit_inR95;
  logic [6:0] lit_inR96;
  logic [6:0] lit_inR97;
  logic [6:0] lit_inR98;
  logic [6:0] lit_inR99;
  logic [6:0] lit_inR100;
  logic [6:0] lit_inR101;
  logic [6:0] lit_inR102;
  logic [6:0] lit_inR103;
  logic [6:0] lit_inR104;
  logic [6:0] lit_inR105;
  logic [6:0] lit_inR106;
  logic [6:0] lit_inR107;
  logic [6:0] lit_inR108;
  logic [6:0] lit_inR109;
  logic [6:0] lit_inR110;
  logic [6:0] lit_inR111;
  logic [6:0] lit_inR112;
  logic [6:0] lit_inR113;
  logic [6:0] lit_inR114;
  logic [6:0] lit_inR115;
  logic [6:0] lit_inR116;
  logic [6:0] lit_inR117;
  logic [6:0] lit_inR118;
  logic [6:0] lit_inR119;
  logic [6:0] lit_inR120;
  logic [6:0] lit_inR121;
  logic [6:0] lit_inR122;
  logic [6:0] lit_inR123;
  logic [6:0] lit_inR124;
  logic [6:0] lit_inR125;
  assign zll_main_nextpc7_in = {arg0, arg0};
  assign zll_main_nextpc5_in = zll_main_nextpc7_in[77:0];
  assign zll_main_nextpc1_in = {zll_main_nextpc5_in[38:0], zll_main_nextpc5_in[77:39]};
  assign zll_main_nextpc3_in = {zll_main_nextpc1_in[38:7], zll_main_nextpc1_in[77:39], zll_main_nextpc1_in[6:0]};
  assign zll_main_nextpc4_in = {zll_main_nextpc3_in[77:46], zll_main_nextpc3_in[6:0], zll_main_nextpc3_in[45:7]};
  assign od19_programcounter_incpc_in = zll_main_nextpc4_in[45:39];
  assign zll_od19_programcounter_incpc213_in = {od19_programcounter_incpc_in[6:0], od19_programcounter_incpc_in[6:0]};
  assign zll_od19_programcounter_incpc129_in = {zll_od19_programcounter_incpc213_in[13:7], zll_od19_programcounter_incpc213_in[13:7]};
  assign zll_od19_programcounter_incpc70_in = {zll_od19_programcounter_incpc129_in[13:7], zll_od19_programcounter_incpc129_in[13:7]};
  assign zll_od19_programcounter_incpc105_in = {zll_od19_programcounter_incpc70_in[13:7], zll_od19_programcounter_incpc70_in[13:7]};
  assign zll_od19_programcounter_incpc2_in = {zll_od19_programcounter_incpc105_in[13:7], zll_od19_programcounter_incpc105_in[13:7]};
  assign zll_od19_programcounter_incpc118_in = {zll_od19_programcounter_incpc2_in[13:7], zll_od19_programcounter_incpc2_in[13:7]};
  assign zll_od19_programcounter_incpc208_in = {zll_od19_programcounter_incpc118_in[13:7], zll_od19_programcounter_incpc118_in[13:7]};
  assign zll_od19_programcounter_incpc172_in = {zll_od19_programcounter_incpc208_in[13:7], zll_od19_programcounter_incpc208_in[13:7]};
  assign zll_od19_programcounter_incpc98_in = {zll_od19_programcounter_incpc172_in[13:7], zll_od19_programcounter_incpc172_in[13:7]};
  assign zll_od19_programcounter_incpc34_in = {zll_od19_programcounter_incpc98_in[13:7], zll_od19_programcounter_incpc98_in[13:7]};
  assign zll_od19_programcounter_incpc116_in = {zll_od19_programcounter_incpc34_in[13:7], zll_od19_programcounter_incpc34_in[13:7]};
  assign zll_od19_programcounter_incpc72_in = {zll_od19_programcounter_incpc116_in[13:7], zll_od19_programcounter_incpc116_in[13:7]};
  assign zll_od19_programcounter_incpc4_in = {zll_od19_programcounter_incpc72_in[13:7], zll_od19_programcounter_incpc72_in[13:7]};
  assign zll_od19_programcounter_incpc148_in = {zll_od19_programcounter_incpc4_in[13:7], zll_od19_programcounter_incpc4_in[13:7]};
  assign zll_od19_programcounter_incpc121_in = {zll_od19_programcounter_incpc148_in[13:7], zll_od19_programcounter_incpc148_in[13:7]};
  assign zll_od19_programcounter_incpc77_in = {zll_od19_programcounter_incpc121_in[13:7], zll_od19_programcounter_incpc121_in[13:7]};
  assign zll_od19_programcounter_incpc12_in = {zll_od19_programcounter_incpc77_in[13:7], zll_od19_programcounter_incpc77_in[13:7]};
  assign zll_od19_programcounter_incpc39_in = {zll_od19_programcounter_incpc12_in[13:7], zll_od19_programcounter_incpc12_in[13:7]};
  assign zll_od19_programcounter_incpc161_in = {zll_od19_programcounter_incpc39_in[13:7], zll_od19_programcounter_incpc39_in[13:7]};
  assign zll_od19_programcounter_incpc26_in = {zll_od19_programcounter_incpc161_in[13:7], zll_od19_programcounter_incpc161_in[13:7]};
  assign zll_od19_programcounter_incpc111_in = {zll_od19_programcounter_incpc26_in[13:7], zll_od19_programcounter_incpc26_in[13:7]};
  assign zll_od19_programcounter_incpc219_in = {zll_od19_programcounter_incpc111_in[13:7], zll_od19_programcounter_incpc111_in[13:7]};
  assign zll_od19_programcounter_incpc8_in = {zll_od19_programcounter_incpc219_in[13:7], zll_od19_programcounter_incpc219_in[13:7]};
  assign zll_od19_programcounter_incpc147_in = {zll_od19_programcounter_incpc8_in[13:7], zll_od19_programcounter_incpc8_in[13:7]};
  assign zll_od19_programcounter_incpc60_in = {zll_od19_programcounter_incpc147_in[13:7], zll_od19_programcounter_incpc147_in[13:7]};
  assign zll_od19_programcounter_incpc202_in = {zll_od19_programcounter_incpc60_in[13:7], zll_od19_programcounter_incpc60_in[13:7]};
  assign zll_od19_programcounter_incpc120_in = {zll_od19_programcounter_incpc202_in[13:7], zll_od19_programcounter_incpc202_in[13:7]};
  assign zll_od19_programcounter_incpc182_in = {zll_od19_programcounter_incpc120_in[13:7], zll_od19_programcounter_incpc120_in[13:7]};
  assign zll_od19_programcounter_incpc114_in = {zll_od19_programcounter_incpc182_in[13:7], zll_od19_programcounter_incpc182_in[13:7]};
  assign zll_od19_programcounter_incpc196_in = {zll_od19_programcounter_incpc114_in[13:7], zll_od19_programcounter_incpc114_in[13:7]};
  assign zll_od19_programcounter_incpc236_in = {zll_od19_programcounter_incpc196_in[13:7], zll_od19_programcounter_incpc196_in[13:7]};
  assign zll_od19_programcounter_incpc164_in = {zll_od19_programcounter_incpc236_in[13:7], zll_od19_programcounter_incpc236_in[13:7]};
  assign zll_od19_programcounter_incpc226_in = {zll_od19_programcounter_incpc164_in[13:7], zll_od19_programcounter_incpc164_in[13:7]};
  assign zll_od19_programcounter_incpc123_in = {zll_od19_programcounter_incpc226_in[13:7], zll_od19_programcounter_incpc226_in[13:7]};
  assign zll_od19_programcounter_incpc55_in = {zll_od19_programcounter_incpc123_in[13:7], zll_od19_programcounter_incpc123_in[13:7]};
  assign zll_od19_programcounter_incpc175_in = {zll_od19_programcounter_incpc55_in[13:7], zll_od19_programcounter_incpc55_in[13:7]};
  assign zll_od19_programcounter_incpc224_in = {zll_od19_programcounter_incpc175_in[13:7], zll_od19_programcounter_incpc175_in[13:7]};
  assign zll_od19_programcounter_incpc71_in = {zll_od19_programcounter_incpc224_in[13:7], zll_od19_programcounter_incpc224_in[13:7]};
  assign zll_od19_programcounter_incpc198_in = {zll_od19_programcounter_incpc71_in[13:7], zll_od19_programcounter_incpc71_in[13:7]};
  assign zll_od19_programcounter_incpc50_in = {zll_od19_programcounter_incpc198_in[13:7], zll_od19_programcounter_incpc198_in[13:7]};
  assign zll_od19_programcounter_incpc128_in = {zll_od19_programcounter_incpc50_in[13:7], zll_od19_programcounter_incpc50_in[13:7]};
  assign zll_od19_programcounter_incpc27_in = {zll_od19_programcounter_incpc128_in[13:7], zll_od19_programcounter_incpc128_in[13:7]};
  assign zll_od19_programcounter_incpc38_in = {zll_od19_programcounter_incpc27_in[13:7], zll_od19_programcounter_incpc27_in[13:7]};
  assign zll_od19_programcounter_incpc173_in = {zll_od19_programcounter_incpc38_in[13:7], zll_od19_programcounter_incpc38_in[13:7]};
  assign zll_od19_programcounter_incpc117_in = {zll_od19_programcounter_incpc173_in[13:7], zll_od19_programcounter_incpc173_in[13:7]};
  assign zll_od19_programcounter_incpc134_in = {zll_od19_programcounter_incpc117_in[13:7], zll_od19_programcounter_incpc117_in[13:7]};
  assign zll_od19_programcounter_incpc59_in = {zll_od19_programcounter_incpc134_in[13:7], zll_od19_programcounter_incpc134_in[13:7]};
  assign zll_od19_programcounter_incpc227_in = {zll_od19_programcounter_incpc59_in[13:7], zll_od19_programcounter_incpc59_in[13:7]};
  assign zll_od19_programcounter_incpc183_in = {zll_od19_programcounter_incpc227_in[13:7], zll_od19_programcounter_incpc227_in[13:7]};
  assign zll_od19_programcounter_incpc253_in = {zll_od19_programcounter_incpc183_in[13:7], zll_od19_programcounter_incpc183_in[13:7]};
  assign zll_od19_programcounter_incpc203_in = {zll_od19_programcounter_incpc253_in[13:7], zll_od19_programcounter_incpc253_in[13:7]};
  assign zll_od19_programcounter_incpc125_in = {zll_od19_programcounter_incpc203_in[13:7], zll_od19_programcounter_incpc203_in[13:7]};
  assign zll_od19_programcounter_incpc144_in = {zll_od19_programcounter_incpc125_in[13:7], zll_od19_programcounter_incpc125_in[13:7]};
  assign zll_od19_programcounter_incpc113_in = {zll_od19_programcounter_incpc144_in[13:7], zll_od19_programcounter_incpc144_in[13:7]};
  assign zll_od19_programcounter_incpc23_in = {zll_od19_programcounter_incpc113_in[13:7], zll_od19_programcounter_incpc113_in[13:7]};
  assign zll_od19_programcounter_incpc231_in = {zll_od19_programcounter_incpc23_in[13:7], zll_od19_programcounter_incpc23_in[13:7]};
  assign zll_od19_programcounter_incpc212_in = {zll_od19_programcounter_incpc231_in[13:7], zll_od19_programcounter_incpc231_in[13:7]};
  assign zll_od19_programcounter_incpc190_in = {zll_od19_programcounter_incpc212_in[13:7], zll_od19_programcounter_incpc212_in[13:7]};
  assign zll_od19_programcounter_incpc245_in = {zll_od19_programcounter_incpc190_in[13:7], zll_od19_programcounter_incpc190_in[13:7]};
  assign zll_od19_programcounter_incpc52_in = {zll_od19_programcounter_incpc245_in[13:7], zll_od19_programcounter_incpc245_in[13:7]};
  assign zll_od19_programcounter_incpc56_in = {zll_od19_programcounter_incpc52_in[13:7], zll_od19_programcounter_incpc52_in[13:7]};
  assign zll_od19_programcounter_incpc131_in = {zll_od19_programcounter_incpc56_in[13:7], zll_od19_programcounter_incpc56_in[13:7]};
  assign zll_od19_programcounter_incpc51_in = {zll_od19_programcounter_incpc131_in[13:7], zll_od19_programcounter_incpc131_in[13:7]};
  assign zll_od19_programcounter_incpc230_in = {zll_od19_programcounter_incpc51_in[13:7], zll_od19_programcounter_incpc51_in[13:7]};
  assign zll_od19_programcounter_incpc168_in = {zll_od19_programcounter_incpc230_in[13:7], zll_od19_programcounter_incpc230_in[13:7]};
  assign zll_od19_programcounter_incpc127_in = {zll_od19_programcounter_incpc168_in[13:7], zll_od19_programcounter_incpc168_in[13:7]};
  assign zll_od19_programcounter_incpc41_in = {zll_od19_programcounter_incpc127_in[13:7], zll_od19_programcounter_incpc127_in[13:7]};
  assign zll_od19_programcounter_incpc18_in = {zll_od19_programcounter_incpc41_in[13:7], zll_od19_programcounter_incpc41_in[13:7]};
  assign zll_od19_programcounter_incpc174_in = {zll_od19_programcounter_incpc18_in[13:7], zll_od19_programcounter_incpc18_in[13:7]};
  assign zll_od19_programcounter_incpc112_in = {zll_od19_programcounter_incpc174_in[13:7], zll_od19_programcounter_incpc174_in[13:7]};
  assign zll_od19_programcounter_incpc24_in = {zll_od19_programcounter_incpc112_in[13:7], zll_od19_programcounter_incpc112_in[13:7]};
  assign zll_od19_programcounter_incpc66_in = {zll_od19_programcounter_incpc24_in[13:7], zll_od19_programcounter_incpc24_in[13:7]};
  assign zll_od19_programcounter_incpc35_in = {zll_od19_programcounter_incpc66_in[13:7], zll_od19_programcounter_incpc66_in[13:7]};
  assign zll_od19_programcounter_incpc215_in = {zll_od19_programcounter_incpc35_in[13:7], zll_od19_programcounter_incpc35_in[13:7]};
  assign zll_od19_programcounter_incpc69_in = {zll_od19_programcounter_incpc215_in[13:7], zll_od19_programcounter_incpc215_in[13:7]};
  assign zll_od19_programcounter_incpc136_in = {zll_od19_programcounter_incpc69_in[13:7], zll_od19_programcounter_incpc69_in[13:7]};
  assign zll_od19_programcounter_incpc187_in = {zll_od19_programcounter_incpc136_in[13:7], zll_od19_programcounter_incpc136_in[13:7]};
  assign zll_od19_programcounter_incpc241_in = {zll_od19_programcounter_incpc187_in[13:7], zll_od19_programcounter_incpc187_in[13:7]};
  assign zll_od19_programcounter_incpc81_in = {zll_od19_programcounter_incpc241_in[13:7], zll_od19_programcounter_incpc241_in[13:7]};
  assign zll_od19_programcounter_incpc169_in = {zll_od19_programcounter_incpc81_in[13:7], zll_od19_programcounter_incpc81_in[13:7]};
  assign zll_od19_programcounter_incpc207_in = {zll_od19_programcounter_incpc169_in[13:7], zll_od19_programcounter_incpc169_in[13:7]};
  assign zll_od19_programcounter_incpc193_in = {zll_od19_programcounter_incpc207_in[13:7], zll_od19_programcounter_incpc207_in[13:7]};
  assign zll_od19_programcounter_incpc218_in = {zll_od19_programcounter_incpc193_in[13:7], zll_od19_programcounter_incpc193_in[13:7]};
  assign zll_od19_programcounter_incpc109_in = {zll_od19_programcounter_incpc218_in[13:7], zll_od19_programcounter_incpc218_in[13:7]};
  assign zll_od19_programcounter_incpc156_in = {zll_od19_programcounter_incpc109_in[13:7], zll_od19_programcounter_incpc109_in[13:7]};
  assign zll_od19_programcounter_incpc115_in = {zll_od19_programcounter_incpc156_in[13:7], zll_od19_programcounter_incpc156_in[13:7]};
  assign zll_od19_programcounter_incpc53_in = {zll_od19_programcounter_incpc115_in[13:7], zll_od19_programcounter_incpc115_in[13:7]};
  assign zll_od19_programcounter_incpc151_in = {zll_od19_programcounter_incpc53_in[13:7], zll_od19_programcounter_incpc53_in[13:7]};
  assign zll_od19_programcounter_incpc63_in = {zll_od19_programcounter_incpc151_in[13:7], zll_od19_programcounter_incpc151_in[13:7]};
  assign zll_od19_programcounter_incpc106_in = {zll_od19_programcounter_incpc63_in[13:7], zll_od19_programcounter_incpc63_in[13:7]};
  assign zll_od19_programcounter_incpc142_in = {zll_od19_programcounter_incpc106_in[13:7], zll_od19_programcounter_incpc106_in[13:7]};
  assign zll_od19_programcounter_incpc191_in = {zll_od19_programcounter_incpc142_in[13:7], zll_od19_programcounter_incpc142_in[13:7]};
  assign zll_od19_programcounter_incpc204_in = {zll_od19_programcounter_incpc191_in[13:7], zll_od19_programcounter_incpc191_in[13:7]};
  assign zll_od19_programcounter_incpc119_in = {zll_od19_programcounter_incpc204_in[13:7], zll_od19_programcounter_incpc204_in[13:7]};
  assign zll_od19_programcounter_incpc90_in = {zll_od19_programcounter_incpc119_in[13:7], zll_od19_programcounter_incpc119_in[13:7]};
  assign zll_od19_programcounter_incpc85_in = {zll_od19_programcounter_incpc90_in[13:7], zll_od19_programcounter_incpc90_in[13:7]};
  assign zll_od19_programcounter_incpc62_in = {zll_od19_programcounter_incpc85_in[13:7], zll_od19_programcounter_incpc85_in[13:7]};
  assign zll_od19_programcounter_incpc94_in = {zll_od19_programcounter_incpc62_in[13:7], zll_od19_programcounter_incpc62_in[13:7]};
  assign zll_od19_programcounter_incpc186_in = {zll_od19_programcounter_incpc94_in[13:7], zll_od19_programcounter_incpc94_in[13:7]};
  assign zll_od19_programcounter_incpc11_in = {zll_od19_programcounter_incpc186_in[13:7], zll_od19_programcounter_incpc186_in[13:7]};
  assign zll_od19_programcounter_incpc37_in = {zll_od19_programcounter_incpc11_in[13:7], zll_od19_programcounter_incpc11_in[13:7]};
  assign zll_od19_programcounter_incpc167_in = {zll_od19_programcounter_incpc37_in[13:7], zll_od19_programcounter_incpc37_in[13:7]};
  assign zll_od19_programcounter_incpc247_in = {zll_od19_programcounter_incpc167_in[13:7], zll_od19_programcounter_incpc167_in[13:7]};
  assign zll_od19_programcounter_incpc185_in = {zll_od19_programcounter_incpc247_in[13:7], zll_od19_programcounter_incpc247_in[13:7]};
  assign zll_od19_programcounter_incpc80_in = {zll_od19_programcounter_incpc185_in[13:7], zll_od19_programcounter_incpc185_in[13:7]};
  assign zll_od19_programcounter_incpc145_in = {zll_od19_programcounter_incpc80_in[13:7], zll_od19_programcounter_incpc80_in[13:7]};
  assign zll_od19_programcounter_incpc10_in = {zll_od19_programcounter_incpc145_in[13:7], zll_od19_programcounter_incpc145_in[13:7]};
  assign zll_od19_programcounter_incpc49_in = {zll_od19_programcounter_incpc10_in[13:7], zll_od19_programcounter_incpc10_in[13:7]};
  assign zll_od19_programcounter_incpc93_in = {zll_od19_programcounter_incpc49_in[13:7], zll_od19_programcounter_incpc49_in[13:7]};
  assign zll_od19_programcounter_incpc91_in = {zll_od19_programcounter_incpc93_in[13:7], zll_od19_programcounter_incpc93_in[13:7]};
  assign zll_od19_programcounter_incpc163_in = {zll_od19_programcounter_incpc91_in[13:7], zll_od19_programcounter_incpc91_in[13:7]};
  assign zll_od19_programcounter_incpc64_in = {zll_od19_programcounter_incpc163_in[13:7], zll_od19_programcounter_incpc163_in[13:7]};
  assign zll_od19_programcounter_incpc101_in = {zll_od19_programcounter_incpc64_in[13:7], zll_od19_programcounter_incpc64_in[13:7]};
  assign zll_od19_programcounter_incpc238_in = {zll_od19_programcounter_incpc101_in[13:7], zll_od19_programcounter_incpc101_in[13:7]};
  assign zll_od19_programcounter_incpc221_in = {zll_od19_programcounter_incpc238_in[13:7], zll_od19_programcounter_incpc238_in[13:7]};
  assign zll_od19_programcounter_incpc78_in = {zll_od19_programcounter_incpc221_in[13:7], zll_od19_programcounter_incpc221_in[13:7]};
  assign zll_od19_programcounter_incpc22_in = {zll_od19_programcounter_incpc78_in[13:7], zll_od19_programcounter_incpc78_in[13:7]};
  assign zll_od19_programcounter_incpc220_in = {zll_od19_programcounter_incpc22_in[13:7], zll_od19_programcounter_incpc22_in[13:7]};
  assign zll_od19_programcounter_incpc97_in = {zll_od19_programcounter_incpc220_in[13:7], zll_od19_programcounter_incpc220_in[13:7]};
  assign zll_od19_programcounter_incpc143_in = {zll_od19_programcounter_incpc97_in[13:7], zll_od19_programcounter_incpc97_in[13:7]};
  assign zll_od19_programcounter_incpc197_in = {zll_od19_programcounter_incpc143_in[13:7], zll_od19_programcounter_incpc143_in[13:7]};
  assign zll_od19_programcounter_incpc194_in = {zll_od19_programcounter_incpc197_in[13:7], zll_od19_programcounter_incpc197_in[13:7]};
  assign zll_od19_programcounter_incpc158_in = {zll_od19_programcounter_incpc194_in[13:7], zll_od19_programcounter_incpc194_in[13:7]};
  assign zll_od19_programcounter_incpc40_in = {zll_od19_programcounter_incpc158_in[13:7], zll_od19_programcounter_incpc158_in[13:7]};
  assign zll_od19_programcounter_incpc250_in = {zll_od19_programcounter_incpc40_in[13:7], zll_od19_programcounter_incpc40_in[13:7]};
  assign zll_od19_programcounter_incpc171_in = {zll_od19_programcounter_incpc250_in[13:7], zll_od19_programcounter_incpc250_in[13:7]};
  assign lit_in = zll_od19_programcounter_incpc171_in[6:0];
  assign lit_inR1 = zll_od19_programcounter_incpc250_in[6:0];
  assign lit_inR2 = zll_od19_programcounter_incpc40_in[6:0];
  assign lit_inR3 = zll_od19_programcounter_incpc158_in[6:0];
  assign lit_inR4 = zll_od19_programcounter_incpc194_in[6:0];
  assign lit_inR5 = zll_od19_programcounter_incpc197_in[6:0];
  assign lit_inR6 = zll_od19_programcounter_incpc143_in[6:0];
  assign lit_inR7 = zll_od19_programcounter_incpc97_in[6:0];
  assign lit_inR8 = zll_od19_programcounter_incpc220_in[6:0];
  assign lit_inR9 = zll_od19_programcounter_incpc22_in[6:0];
  assign lit_inR10 = zll_od19_programcounter_incpc78_in[6:0];
  assign lit_inR11 = zll_od19_programcounter_incpc221_in[6:0];
  assign lit_inR12 = zll_od19_programcounter_incpc238_in[6:0];
  assign lit_inR13 = zll_od19_programcounter_incpc101_in[6:0];
  assign lit_inR14 = zll_od19_programcounter_incpc64_in[6:0];
  assign lit_inR15 = zll_od19_programcounter_incpc163_in[6:0];
  assign lit_inR16 = zll_od19_programcounter_incpc91_in[6:0];
  assign lit_inR17 = zll_od19_programcounter_incpc93_in[6:0];
  assign lit_inR18 = zll_od19_programcounter_incpc49_in[6:0];
  assign lit_inR19 = zll_od19_programcounter_incpc10_in[6:0];
  assign lit_inR20 = zll_od19_programcounter_incpc145_in[6:0];
  assign lit_inR21 = zll_od19_programcounter_incpc80_in[6:0];
  assign lit_inR22 = zll_od19_programcounter_incpc185_in[6:0];
  assign lit_inR23 = zll_od19_programcounter_incpc247_in[6:0];
  assign lit_inR24 = zll_od19_programcounter_incpc167_in[6:0];
  assign lit_inR25 = zll_od19_programcounter_incpc37_in[6:0];
  assign lit_inR26 = zll_od19_programcounter_incpc11_in[6:0];
  assign lit_inR27 = zll_od19_programcounter_incpc186_in[6:0];
  assign lit_inR28 = zll_od19_programcounter_incpc94_in[6:0];
  assign lit_inR29 = zll_od19_programcounter_incpc62_in[6:0];
  assign lit_inR30 = zll_od19_programcounter_incpc85_in[6:0];
  assign lit_inR31 = zll_od19_programcounter_incpc90_in[6:0];
  assign lit_inR32 = zll_od19_programcounter_incpc119_in[6:0];
  assign lit_inR33 = zll_od19_programcounter_incpc204_in[6:0];
  assign lit_inR34 = zll_od19_programcounter_incpc191_in[6:0];
  assign lit_inR35 = zll_od19_programcounter_incpc142_in[6:0];
  assign lit_inR36 = zll_od19_programcounter_incpc106_in[6:0];
  assign lit_inR37 = zll_od19_programcounter_incpc63_in[6:0];
  assign lit_inR38 = zll_od19_programcounter_incpc151_in[6:0];
  assign lit_inR39 = zll_od19_programcounter_incpc53_in[6:0];
  assign lit_inR40 = zll_od19_programcounter_incpc115_in[6:0];
  assign lit_inR41 = zll_od19_programcounter_incpc156_in[6:0];
  assign lit_inR42 = zll_od19_programcounter_incpc109_in[6:0];
  assign lit_inR43 = zll_od19_programcounter_incpc218_in[6:0];
  assign lit_inR44 = zll_od19_programcounter_incpc193_in[6:0];
  assign lit_inR45 = zll_od19_programcounter_incpc207_in[6:0];
  assign lit_inR46 = zll_od19_programcounter_incpc169_in[6:0];
  assign lit_inR47 = zll_od19_programcounter_incpc81_in[6:0];
  assign lit_inR48 = zll_od19_programcounter_incpc241_in[6:0];
  assign lit_inR49 = zll_od19_programcounter_incpc187_in[6:0];
  assign lit_inR50 = zll_od19_programcounter_incpc136_in[6:0];
  assign lit_inR51 = zll_od19_programcounter_incpc69_in[6:0];
  assign lit_inR52 = zll_od19_programcounter_incpc215_in[6:0];
  assign lit_inR53 = zll_od19_programcounter_incpc35_in[6:0];
  assign lit_inR54 = zll_od19_programcounter_incpc66_in[6:0];
  assign lit_inR55 = zll_od19_programcounter_incpc24_in[6:0];
  assign lit_inR56 = zll_od19_programcounter_incpc112_in[6:0];
  assign lit_inR57 = zll_od19_programcounter_incpc174_in[6:0];
  assign lit_inR58 = zll_od19_programcounter_incpc18_in[6:0];
  assign lit_inR59 = zll_od19_programcounter_incpc41_in[6:0];
  assign lit_inR60 = zll_od19_programcounter_incpc127_in[6:0];
  assign lit_inR61 = zll_od19_programcounter_incpc168_in[6:0];
  assign lit_inR62 = zll_od19_programcounter_incpc230_in[6:0];
  assign lit_inR63 = zll_od19_programcounter_incpc51_in[6:0];
  assign lit_inR64 = zll_od19_programcounter_incpc131_in[6:0];
  assign lit_inR65 = zll_od19_programcounter_incpc56_in[6:0];
  assign lit_inR66 = zll_od19_programcounter_incpc52_in[6:0];
  assign lit_inR67 = zll_od19_programcounter_incpc245_in[6:0];
  assign lit_inR68 = zll_od19_programcounter_incpc190_in[6:0];
  assign lit_inR69 = zll_od19_programcounter_incpc212_in[6:0];
  assign lit_inR70 = zll_od19_programcounter_incpc231_in[6:0];
  assign lit_inR71 = zll_od19_programcounter_incpc23_in[6:0];
  assign lit_inR72 = zll_od19_programcounter_incpc113_in[6:0];
  assign lit_inR73 = zll_od19_programcounter_incpc144_in[6:0];
  assign lit_inR74 = zll_od19_programcounter_incpc125_in[6:0];
  assign lit_inR75 = zll_od19_programcounter_incpc203_in[6:0];
  assign lit_inR76 = zll_od19_programcounter_incpc253_in[6:0];
  assign lit_inR77 = zll_od19_programcounter_incpc183_in[6:0];
  assign lit_inR78 = zll_od19_programcounter_incpc227_in[6:0];
  assign lit_inR79 = zll_od19_programcounter_incpc59_in[6:0];
  assign lit_inR80 = zll_od19_programcounter_incpc134_in[6:0];
  assign lit_inR81 = zll_od19_programcounter_incpc117_in[6:0];
  assign lit_inR82 = zll_od19_programcounter_incpc173_in[6:0];
  assign lit_inR83 = zll_od19_programcounter_incpc38_in[6:0];
  assign lit_inR84 = zll_od19_programcounter_incpc27_in[6:0];
  assign lit_inR85 = zll_od19_programcounter_incpc128_in[6:0];
  assign lit_inR86 = zll_od19_programcounter_incpc50_in[6:0];
  assign lit_inR87 = zll_od19_programcounter_incpc198_in[6:0];
  assign lit_inR88 = zll_od19_programcounter_incpc71_in[6:0];
  assign lit_inR89 = zll_od19_programcounter_incpc224_in[6:0];
  assign lit_inR90 = zll_od19_programcounter_incpc175_in[6:0];
  assign lit_inR91 = zll_od19_programcounter_incpc55_in[6:0];
  assign lit_inR92 = zll_od19_programcounter_incpc123_in[6:0];
  assign lit_inR93 = zll_od19_programcounter_incpc226_in[6:0];
  assign lit_inR94 = zll_od19_programcounter_incpc164_in[6:0];
  assign lit_inR95 = zll_od19_programcounter_incpc236_in[6:0];
  assign lit_inR96 = zll_od19_programcounter_incpc196_in[6:0];
  assign lit_inR97 = zll_od19_programcounter_incpc114_in[6:0];
  assign lit_inR98 = zll_od19_programcounter_incpc182_in[6:0];
  assign lit_inR99 = zll_od19_programcounter_incpc120_in[6:0];
  assign lit_inR100 = zll_od19_programcounter_incpc202_in[6:0];
  assign lit_inR101 = zll_od19_programcounter_incpc60_in[6:0];
  assign lit_inR102 = zll_od19_programcounter_incpc147_in[6:0];
  assign lit_inR103 = zll_od19_programcounter_incpc8_in[6:0];
  assign lit_inR104 = zll_od19_programcounter_incpc219_in[6:0];
  assign lit_inR105 = zll_od19_programcounter_incpc111_in[6:0];
  assign lit_inR106 = zll_od19_programcounter_incpc26_in[6:0];
  assign lit_inR107 = zll_od19_programcounter_incpc161_in[6:0];
  assign lit_inR108 = zll_od19_programcounter_incpc39_in[6:0];
  assign lit_inR109 = zll_od19_programcounter_incpc12_in[6:0];
  assign lit_inR110 = zll_od19_programcounter_incpc77_in[6:0];
  assign lit_inR111 = zll_od19_programcounter_incpc121_in[6:0];
  assign lit_inR112 = zll_od19_programcounter_incpc148_in[6:0];
  assign lit_inR113 = zll_od19_programcounter_incpc4_in[6:0];
  assign lit_inR114 = zll_od19_programcounter_incpc72_in[6:0];
  assign lit_inR115 = zll_od19_programcounter_incpc116_in[6:0];
  assign lit_inR116 = zll_od19_programcounter_incpc34_in[6:0];
  assign lit_inR117 = zll_od19_programcounter_incpc98_in[6:0];
  assign lit_inR118 = zll_od19_programcounter_incpc172_in[6:0];
  assign lit_inR119 = zll_od19_programcounter_incpc208_in[6:0];
  assign lit_inR120 = zll_od19_programcounter_incpc118_in[6:0];
  assign lit_inR121 = zll_od19_programcounter_incpc2_in[6:0];
  assign lit_inR122 = zll_od19_programcounter_incpc105_in[6:0];
  assign lit_inR123 = zll_od19_programcounter_incpc70_in[6:0];
  assign lit_inR124 = zll_od19_programcounter_incpc129_in[6:0];
  assign lit_inR125 = zll_od19_programcounter_incpc213_in[6:0];
  assign res = {zll_main_nextpc4_in[77:46], (lit_inR125[6:0] == 7'h0) ? 7'h1 : ((lit_inR124[6:0] == 7'h1) ? 7'h2 : ((lit_inR123[6:0] == 7'h2) ? 7'h3 : ((lit_inR122[6:0] == 7'h3) ? 7'h4 : ((lit_inR121[6:0] == 7'h4) ? 7'h5 : ((lit_inR120[6:0] == 7'h5) ? 7'h6 : ((lit_inR119[6:0] == 7'h6) ? 7'h7 : ((lit_inR118[6:0] == 7'h7) ? 7'h8 : ((lit_inR117[6:0] == 7'h8) ? 7'h9 : ((lit_inR116[6:0] == 7'h9) ? 7'ha : ((lit_inR115[6:0] == 7'ha) ? 7'hb : ((lit_inR114[6:0] == 7'hb) ? 7'hc : ((lit_inR113[6:0] == 7'hc) ? 7'hd : ((lit_inR112[6:0] == 7'hd) ? 7'he : ((lit_inR111[6:0] == 7'he) ? 7'hf : ((lit_inR110[6:0] == 7'hf) ? 7'h10 : ((lit_inR109[6:0] == 7'h10) ? 7'h11 : ((lit_inR108[6:0] == 7'h11) ? 7'h12 : ((lit_inR107[6:0] == 7'h12) ? 7'h13 : ((lit_inR106[6:0] == 7'h13) ? 7'h14 : ((lit_inR105[6:0] == 7'h14) ? 7'h15 : ((lit_inR104[6:0] == 7'h15) ? 7'h16 : ((lit_inR103[6:0] == 7'h16) ? 7'h17 : ((lit_inR102[6:0] == 7'h17) ? 7'h18 : ((lit_inR101[6:0] == 7'h18) ? 7'h19 : ((lit_inR100[6:0] == 7'h19) ? 7'h1a : ((lit_inR99[6:0] == 7'h1a) ? 7'h1b : ((lit_inR98[6:0] == 7'h1b) ? 7'h1c : ((lit_inR97[6:0] == 7'h1c) ? 7'h1d : ((lit_inR96[6:0] == 7'h1d) ? 7'h1e : ((lit_inR95[6:0] == 7'h1e) ? 7'h1f : ((lit_inR94[6:0] == 7'h1f) ? 7'h20 : ((lit_inR93[6:0] == 7'h20) ? 7'h21 : ((lit_inR92[6:0] == 7'h21) ? 7'h22 : ((lit_inR91[6:0] == 7'h22) ? 7'h23 : ((lit_inR90[6:0] == 7'h23) ? 7'h24 : ((lit_inR89[6:0] == 7'h24) ? 7'h25 : ((lit_inR88[6:0] == 7'h25) ? 7'h26 : ((lit_inR87[6:0] == 7'h26) ? 7'h27 : ((lit_inR86[6:0] == 7'h27) ? 7'h28 : ((lit_inR85[6:0] == 7'h28) ? 7'h29 : ((lit_inR84[6:0] == 7'h29) ? 7'h2a : ((lit_inR83[6:0] == 7'h2a) ? 7'h2b : ((lit_inR82[6:0] == 7'h2b) ? 7'h2c : ((lit_inR81[6:0] == 7'h2c) ? 7'h2d : ((lit_inR80[6:0] == 7'h2d) ? 7'h2e : ((lit_inR79[6:0] == 7'h2e) ? 7'h2f : ((lit_inR78[6:0] == 7'h2f) ? 7'h30 : ((lit_inR77[6:0] == 7'h30) ? 7'h31 : ((lit_inR76[6:0] == 7'h31) ? 7'h32 : ((lit_inR75[6:0] == 7'h32) ? 7'h33 : ((lit_inR74[6:0] == 7'h33) ? 7'h34 : ((lit_inR73[6:0] == 7'h34) ? 7'h35 : ((lit_inR72[6:0] == 7'h35) ? 7'h36 : ((lit_inR71[6:0] == 7'h36) ? 7'h37 : ((lit_inR70[6:0] == 7'h37) ? 7'h38 : ((lit_inR69[6:0] == 7'h38) ? 7'h39 : ((lit_inR68[6:0] == 7'h39) ? 7'h3a : ((lit_inR67[6:0] == 7'h3a) ? 7'h3b : ((lit_inR66[6:0] == 7'h3b) ? 7'h3c : ((lit_inR65[6:0] == 7'h3c) ? 7'h3d : ((lit_inR64[6:0] == 7'h3d) ? 7'h3e : ((lit_inR63[6:0] == 7'h3e) ? 7'h3f : ((lit_inR62[6:0] == 7'h3f) ? 7'h40 : ((lit_inR61[6:0] == 7'h40) ? 7'h41 : ((lit_inR60[6:0] == 7'h41) ? 7'h42 : ((lit_inR59[6:0] == 7'h42) ? 7'h43 : ((lit_inR58[6:0] == 7'h43) ? 7'h44 : ((lit_inR57[6:0] == 7'h44) ? 7'h45 : ((lit_inR56[6:0] == 7'h45) ? 7'h46 : ((lit_inR55[6:0] == 7'h46) ? 7'h47 : ((lit_inR54[6:0] == 7'h47) ? 7'h48 : ((lit_inR53[6:0] == 7'h48) ? 7'h49 : ((lit_inR52[6:0] == 7'h49) ? 7'h4a : ((lit_inR51[6:0] == 7'h4a) ? 7'h4b : ((lit_inR50[6:0] == 7'h4b) ? 7'h4c : ((lit_inR49[6:0] == 7'h4c) ? 7'h4d : ((lit_inR48[6:0] == 7'h4d) ? 7'h4e : ((lit_inR47[6:0] == 7'h4e) ? 7'h4f : ((lit_inR46[6:0] == 7'h4f) ? 7'h50 : ((lit_inR45[6:0] == 7'h50) ? 7'h51 : ((lit_inR44[6:0] == 7'h51) ? 7'h52 : ((lit_inR43[6:0] == 7'h52) ? 7'h53 : ((lit_inR42[6:0] == 7'h53) ? 7'h54 : ((lit_inR41[6:0] == 7'h54) ? 7'h55 : ((lit_inR40[6:0] == 7'h55) ? 7'h56 : ((lit_inR39[6:0] == 7'h56) ? 7'h57 : ((lit_inR38[6:0] == 7'h57) ? 7'h58 : ((lit_inR37[6:0] == 7'h58) ? 7'h59 : ((lit_inR36[6:0] == 7'h59) ? 7'h5a : ((lit_inR35[6:0] == 7'h5a) ? 7'h5b : ((lit_inR34[6:0] == 7'h5b) ? 7'h5c : ((lit_inR33[6:0] == 7'h5c) ? 7'h5d : ((lit_inR32[6:0] == 7'h5d) ? 7'h5e : ((lit_inR31[6:0] == 7'h5e) ? 7'h5f : ((lit_inR30[6:0] == 7'h5f) ? 7'h60 : ((lit_inR29[6:0] == 7'h60) ? 7'h61 : ((lit_inR28[6:0] == 7'h61) ? 7'h62 : ((lit_inR27[6:0] == 7'h62) ? 7'h63 : ((lit_inR26[6:0] == 7'h63) ? 7'h64 : ((lit_inR25[6:0] == 7'h64) ? 7'h65 : ((lit_inR24[6:0] == 7'h65) ? 7'h66 : ((lit_inR23[6:0] == 7'h66) ? 7'h67 : ((lit_inR22[6:0] == 7'h67) ? 7'h68 : ((lit_inR21[6:0] == 7'h68) ? 7'h69 : ((lit_inR20[6:0] == 7'h69) ? 7'h6a : ((lit_inR19[6:0] == 7'h6a) ? 7'h6b : ((lit_inR18[6:0] == 7'h6b) ? 7'h6c : ((lit_inR17[6:0] == 7'h6c) ? 7'h6d : ((lit_inR16[6:0] == 7'h6d) ? 7'h6e : ((lit_inR15[6:0] == 7'h6e) ? 7'h6f : ((lit_inR14[6:0] == 7'h6f) ? 7'h70 : ((lit_inR13[6:0] == 7'h70) ? 7'h71 : ((lit_inR12[6:0] == 7'h71) ? 7'h72 : ((lit_inR11[6:0] == 7'h72) ? 7'h73 : ((lit_inR10[6:0] == 7'h73) ? 7'h74 : ((lit_inR9[6:0] == 7'h74) ? 7'h75 : ((lit_inR8[6:0] == 7'h75) ? 7'h76 : ((lit_inR7[6:0] == 7'h76) ? 7'h77 : ((lit_inR6[6:0] == 7'h77) ? 7'h78 : ((lit_inR5[6:0] == 7'h78) ? 7'h79 : ((lit_inR4[6:0] == 7'h79) ? 7'h7a : ((lit_inR3[6:0] == 7'h7a) ? 7'h7b : ((lit_inR2[6:0] == 7'h7b) ? 7'h7c : ((lit_inR1[6:0] == 7'h7c) ? 7'h7d : ((lit_in[6:0] == 7'h7d) ? 7'h7e : 7'h0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))};
endmodule