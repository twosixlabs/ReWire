module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [63:0] __in0,
  input logic [63:0] __in1,
  output logic [63:0] __out0,
  output logic [63:0] __out1);
  logic [127:0] gMainziloop;
  logic [127:0] gMainzicompute;
  logic [127:0] gzdLLziMainzicompute42;
  logic [130:0] gzdLLziMainzicompute20;
  logic [7:0] callRes;
  logic [130:0] gzdLLziMainzicompute20R1;
  logic [7:0] callResR1;
  logic [130:0] gzdLLziMainzicompute20R2;
  logic [7:0] callResR2;
  logic [130:0] gzdLLziMainzicompute20R3;
  logic [7:0] callResR3;
  logic [130:0] gzdLLziMainzicompute20R4;
  logic [7:0] callResR4;
  logic [130:0] gzdLLziMainzicompute20R5;
  logic [7:0] callResR5;
  logic [130:0] gzdLLziMainzicompute20R6;
  logic [7:0] callResR6;
  logic [130:0] gzdLLziMainzicompute20R7;
  logic [7:0] callResR7;
  logic [130:0] gzdLLziMainzicompute41;
  logic [7:0] callResR8;
  logic [130:0] gzdLLziMainzicompute41R1;
  logic [7:0] callResR9;
  logic [130:0] gzdLLziMainzicompute41R2;
  logic [7:0] callResR10;
  logic [130:0] gzdLLziMainzicompute41R3;
  logic [7:0] callResR11;
  logic [130:0] gzdLLziMainzicompute41R4;
  logic [7:0] callResR12;
  logic [130:0] gzdLLziMainzicompute41R5;
  logic [7:0] callResR13;
  logic [130:0] gzdLLziMainzicompute41R6;
  logic [7:0] callResR14;
  logic [130:0] gzdLLziMainzicompute41R7;
  logic [7:0] callResR15;
  logic [128:0] gzdLLziMainziloop2;
  logic [128:0] gzdLLziMainziloop;
  logic [0:0] __continue;
  logic [127:0] __resumption_tag;
  logic [127:0] __resumption_tag_next;
  assign gMainziloop = __resumption_tag;
  assign gMainzicompute = gMainziloop[127:0];
  assign gzdLLziMainzicompute42 = gMainzicompute[127:0];
  assign gzdLLziMainzicompute20 = {gzdLLziMainzicompute42[127:64], gzdLLziMainzicompute42[63:0], 3'h0};
  zdLLziMainzicompute20  zdLLziMainzicompute20 (gzdLLziMainzicompute20[130:67], gzdLLziMainzicompute20[66:3], gzdLLziMainzicompute20[2:0], callRes);
  assign gzdLLziMainzicompute20R1 = {gzdLLziMainzicompute42[127:64], gzdLLziMainzicompute42[63:0], 3'h1};
  zdLLziMainzicompute20  zdLLziMainzicompute20R1 (gzdLLziMainzicompute20R1[130:67], gzdLLziMainzicompute20R1[66:3], gzdLLziMainzicompute20R1[2:0], callResR1);
  assign gzdLLziMainzicompute20R2 = {gzdLLziMainzicompute42[127:64], gzdLLziMainzicompute42[63:0], 3'h2};
  zdLLziMainzicompute20  zdLLziMainzicompute20R2 (gzdLLziMainzicompute20R2[130:67], gzdLLziMainzicompute20R2[66:3], gzdLLziMainzicompute20R2[2:0], callResR2);
  assign gzdLLziMainzicompute20R3 = {gzdLLziMainzicompute42[127:64], gzdLLziMainzicompute42[63:0], 3'h3};
  zdLLziMainzicompute20  zdLLziMainzicompute20R3 (gzdLLziMainzicompute20R3[130:67], gzdLLziMainzicompute20R3[66:3], gzdLLziMainzicompute20R3[2:0], callResR3);
  assign gzdLLziMainzicompute20R4 = {gzdLLziMainzicompute42[127:64], gzdLLziMainzicompute42[63:0], 3'h4};
  zdLLziMainzicompute20  zdLLziMainzicompute20R4 (gzdLLziMainzicompute20R4[130:67], gzdLLziMainzicompute20R4[66:3], gzdLLziMainzicompute20R4[2:0], callResR4);
  assign gzdLLziMainzicompute20R5 = {gzdLLziMainzicompute42[127:64], gzdLLziMainzicompute42[63:0], 3'h5};
  zdLLziMainzicompute20  zdLLziMainzicompute20R5 (gzdLLziMainzicompute20R5[130:67], gzdLLziMainzicompute20R5[66:3], gzdLLziMainzicompute20R5[2:0], callResR5);
  assign gzdLLziMainzicompute20R6 = {gzdLLziMainzicompute42[127:64], gzdLLziMainzicompute42[63:0], 3'h6};
  zdLLziMainzicompute20  zdLLziMainzicompute20R6 (gzdLLziMainzicompute20R6[130:67], gzdLLziMainzicompute20R6[66:3], gzdLLziMainzicompute20R6[2:0], callResR6);
  assign gzdLLziMainzicompute20R7 = {gzdLLziMainzicompute42[127:64], gzdLLziMainzicompute42[63:0], 3'h7};
  zdLLziMainzicompute20  zdLLziMainzicompute20R7 (gzdLLziMainzicompute20R7[130:67], gzdLLziMainzicompute20R7[66:3], gzdLLziMainzicompute20R7[2:0], callResR7);
  assign gzdLLziMainzicompute41 = {gzdLLziMainzicompute42[127:64], gzdLLziMainzicompute42[63:0], 3'h0};
  zdLLziMainzicompute41  zdLLziMainzicompute41 (gzdLLziMainzicompute41[130:67], gzdLLziMainzicompute41[66:3], gzdLLziMainzicompute41[2:0], callResR8);
  assign gzdLLziMainzicompute41R1 = {gzdLLziMainzicompute42[127:64], gzdLLziMainzicompute42[63:0], 3'h1};
  zdLLziMainzicompute41  zdLLziMainzicompute41R1 (gzdLLziMainzicompute41R1[130:67], gzdLLziMainzicompute41R1[66:3], gzdLLziMainzicompute41R1[2:0], callResR9);
  assign gzdLLziMainzicompute41R2 = {gzdLLziMainzicompute42[127:64], gzdLLziMainzicompute42[63:0], 3'h2};
  zdLLziMainzicompute41  zdLLziMainzicompute41R2 (gzdLLziMainzicompute41R2[130:67], gzdLLziMainzicompute41R2[66:3], gzdLLziMainzicompute41R2[2:0], callResR10);
  assign gzdLLziMainzicompute41R3 = {gzdLLziMainzicompute42[127:64], gzdLLziMainzicompute42[63:0], 3'h3};
  zdLLziMainzicompute41  zdLLziMainzicompute41R3 (gzdLLziMainzicompute41R3[130:67], gzdLLziMainzicompute41R3[66:3], gzdLLziMainzicompute41R3[2:0], callResR11);
  assign gzdLLziMainzicompute41R4 = {gzdLLziMainzicompute42[127:64], gzdLLziMainzicompute42[63:0], 3'h4};
  zdLLziMainzicompute41  zdLLziMainzicompute41R4 (gzdLLziMainzicompute41R4[130:67], gzdLLziMainzicompute41R4[66:3], gzdLLziMainzicompute41R4[2:0], callResR12);
  assign gzdLLziMainzicompute41R5 = {gzdLLziMainzicompute42[127:64], gzdLLziMainzicompute42[63:0], 3'h5};
  zdLLziMainzicompute41  zdLLziMainzicompute41R5 (gzdLLziMainzicompute41R5[130:67], gzdLLziMainzicompute41R5[66:3], gzdLLziMainzicompute41R5[2:0], callResR13);
  assign gzdLLziMainzicompute41R6 = {gzdLLziMainzicompute42[127:64], gzdLLziMainzicompute42[63:0], 3'h6};
  zdLLziMainzicompute41  zdLLziMainzicompute41R6 (gzdLLziMainzicompute41R6[130:67], gzdLLziMainzicompute41R6[66:3], gzdLLziMainzicompute41R6[2:0], callResR14);
  assign gzdLLziMainzicompute41R7 = {gzdLLziMainzicompute42[127:64], gzdLLziMainzicompute42[63:0], 3'h7};
  zdLLziMainzicompute41  zdLLziMainzicompute41R7 (gzdLLziMainzicompute41R7[130:67], gzdLLziMainzicompute41R7[66:3], gzdLLziMainzicompute41R7[2:0], callResR15);
  assign gzdLLziMainziloop2 = {1'h0, {callRes, callResR1, callResR2, callResR3, callResR4, callResR5, callResR6, callResR7, callResR8, callResR9, callResR10, callResR11, callResR12, callResR13, callResR14, callResR15}};
  assign gzdLLziMainziloop = gzdLLziMainziloop2[128:0];
  assign {__continue, __out0, __out1, __resumption_tag_next} = {1'h1, gzdLLziMainziloop[127:0]};
  initial __resumption_tag <= {8'h80{1'h0}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      __resumption_tag <= {8'h80{1'h0}};
    end else begin
      __resumption_tag <= __resumption_tag_next;
    end
  end
endmodule

module zdLLziMainzicompute (input logic [63:0] arg0,
  input logic [2:0] arg1,
  output logic [7:0] res);
  logic [63:0] resizze;
  logic [2:0] resizzeR1;
  logic [255:0] binOp;
  logic [255:0] binOpR1;
  logic [127:0] resizzeR2;
  logic [2:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [127:0] resizzeR6;
  assign resizze = arg0;
  assign resizzeR1 = arg1;
  assign binOp = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR1 = {binOp[255:128] * binOp[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR2 = binOpR1[255:128] % binOpR1[127:0];
  assign resizzeR3 = resizzeR2[2:0];
  assign binOpR2 = {128'(resizzeR3[2:0]), 128'h00000000000000000000000000000001};
  assign binOpR3 = {binOpR2[255:128] + binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[2:0];
  assign binOpR4 = {128'h00000000000000000000000000000008, 128'(resizzeR5[2:0])};
  assign binOpR5 = {binOpR4[255:128] - binOpR4[127:0], 128'h00000000000000000000000000000001};
  assign binOpR6 = {binOpR5[255:128] - binOpR5[127:0], 128'h00000000000000000000000000000008};
  assign binOpR7 = {128'(resizze[63:0]), binOpR6[255:128] * binOpR6[127:0]};
  assign resizzeR6 = binOpR7[255:128] >> binOpR7[127:0];
  assign res = resizzeR6[7:0];
endmodule

module zdLLziMainzicompute1 (input logic [63:0] arg0,
  input logic [2:0] arg1,
  output logic [7:0] res);
  logic [63:0] resizze;
  logic [2:0] resizzeR1;
  logic [255:0] binOp;
  logic [255:0] binOpR1;
  logic [127:0] resizzeR2;
  logic [2:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR6;
  logic [2:0] resizzeR7;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [127:0] resizzeR8;
  assign resizze = arg0;
  assign resizzeR1 = arg1;
  assign binOp = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign binOpR1 = {binOp[255:128] - binOp[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR2 = binOpR1[255:128] % binOpR1[127:0];
  assign resizzeR3 = resizzeR2[2:0];
  assign binOpR2 = {128'(resizzeR3[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR3 = {binOpR2[255:128] * binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[2:0];
  assign binOpR4 = {128'(resizzeR5[2:0]), 128'h00000000000000000000000000000001};
  assign binOpR5 = {binOpR4[255:128] + binOpR4[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR6 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR7 = resizzeR6[2:0];
  assign binOpR6 = {128'h00000000000000000000000000000008, 128'(resizzeR7[2:0])};
  assign binOpR7 = {binOpR6[255:128] - binOpR6[127:0], 128'h00000000000000000000000000000001};
  assign binOpR8 = {binOpR7[255:128] - binOpR7[127:0], 128'h00000000000000000000000000000008};
  assign binOpR9 = {128'(resizze[63:0]), binOpR8[255:128] * binOpR8[127:0]};
  assign resizzeR8 = binOpR9[255:128] >> binOpR9[127:0];
  assign res = resizzeR8[7:0];
endmodule

module zdLLziMainzicompute2 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [67:0] gzdLLziMainzicompute1;
  logic [7:0] callRes;
  logic [67:0] gzdLLziMainzicompute;
  logic [7:0] callResR1;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLziMainzicompute1 = {arg1, arg2, binOpR1[255:128] < binOpR1[127:0]};
  zdLLziMainzicompute1  zdLLziMainzicompute1 (gzdLLziMainzicompute1[67:4], gzdLLziMainzicompute1[3:1], callRes);
  assign gzdLLziMainzicompute = {arg0, arg2, binOp[255:128] < binOp[127:0]};
  zdLLziMainzicompute  zdLLziMainzicompute (gzdLLziMainzicompute[67:4], gzdLLziMainzicompute[3:1], callResR1);
  assign res = (gzdLLziMainzicompute[0] == 1'h1) ? callResR1 : callRes;
endmodule

module zdLLziMainzicompute6 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [67:0] gzdLLziMainzicompute5;
  logic [63:0] resizzeR2;
  logic [2:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR6;
  logic [2:0] resizzeR7;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [127:0] resizzeR8;
  logic [67:0] gzdLLziMainzicompute4;
  logic [63:0] resizzeR9;
  logic [2:0] resizzeR10;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [127:0] resizzeR11;
  logic [2:0] resizzeR12;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [255:0] binOpR14;
  logic [255:0] binOpR15;
  logic [127:0] resizzeR13;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLziMainzicompute5 = {arg2, arg1, binOpR1[255:128] < binOpR1[127:0]};
  assign resizzeR2 = gzdLLziMainzicompute5[64:1];
  assign resizzeR3 = gzdLLziMainzicompute5[67:65];
  assign binOpR2 = {128'(resizzeR3[2:0]), 128'h00000000000000000000000000000003};
  assign binOpR3 = {binOpR2[255:128] - binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[2:0];
  assign binOpR4 = {128'(resizzeR5[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR5 = {binOpR4[255:128] * binOpR4[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR6 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR7 = resizzeR6[2:0];
  assign binOpR6 = {128'h00000000000000000000000000000008, 128'(resizzeR7[2:0])};
  assign binOpR7 = {binOpR6[255:128] - binOpR6[127:0], 128'h00000000000000000000000000000001};
  assign binOpR8 = {binOpR7[255:128] - binOpR7[127:0], 128'h00000000000000000000000000000008};
  assign binOpR9 = {128'(resizzeR2[63:0]), binOpR8[255:128] * binOpR8[127:0]};
  assign resizzeR8 = binOpR9[255:128] >> binOpR9[127:0];
  assign gzdLLziMainzicompute4 = {arg2, arg0, binOp[255:128] < binOp[127:0]};
  assign resizzeR9 = gzdLLziMainzicompute4[64:1];
  assign resizzeR10 = gzdLLziMainzicompute4[67:65];
  assign binOpR10 = {128'(resizzeR10[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR11 = {binOpR10[255:128] * binOpR10[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR11 = binOpR11[255:128] % binOpR11[127:0];
  assign resizzeR12 = resizzeR11[2:0];
  assign binOpR12 = {128'h00000000000000000000000000000008, 128'(resizzeR12[2:0])};
  assign binOpR13 = {binOpR12[255:128] - binOpR12[127:0], 128'h00000000000000000000000000000001};
  assign binOpR14 = {binOpR13[255:128] - binOpR13[127:0], 128'h00000000000000000000000000000008};
  assign binOpR15 = {128'(resizzeR9[63:0]), binOpR14[255:128] * binOpR14[127:0]};
  assign resizzeR13 = binOpR15[255:128] >> binOpR15[127:0];
  assign res = (gzdLLziMainzicompute4[0] == 1'h1) ? resizzeR13[7:0] : resizzeR8[7:0];
endmodule

module zdLLziMainzicompute8 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [131:0] gzdLLziMainzicompute7;
  logic [130:0] gzdLLziMainzicompute6;
  logic [7:0] callRes;
  logic [130:0] gzdLLziMainzicompute6R1;
  logic [7:0] callResR1;
  logic [130:0] gzdLLziMainzicompute6R2;
  logic [7:0] callResR2;
  logic [130:0] gzdLLziMainzicompute6R3;
  logic [7:0] callResR3;
  logic [130:0] gzdLLziMainzicompute6R4;
  logic [7:0] callResR4;
  logic [130:0] gzdLLziMainzicompute6R5;
  logic [7:0] callResR5;
  logic [130:0] gzdLLziMainzicompute6R6;
  logic [7:0] callResR6;
  logic [130:0] gzdLLziMainzicompute6R7;
  logic [7:0] callResR7;
  logic [63:0] resizzeR2;
  logic [2:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR6;
  logic [2:0] resizzeR7;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [127:0] resizzeR8;
  logic [131:0] gzdLLziMainzicompute3;
  logic [130:0] gzdLLziMainzicompute2;
  logic [7:0] callResR8;
  logic [130:0] gzdLLziMainzicompute2R1;
  logic [7:0] callResR9;
  logic [130:0] gzdLLziMainzicompute2R2;
  logic [7:0] callResR10;
  logic [130:0] gzdLLziMainzicompute2R3;
  logic [7:0] callResR11;
  logic [130:0] gzdLLziMainzicompute2R4;
  logic [7:0] callResR12;
  logic [130:0] gzdLLziMainzicompute2R5;
  logic [7:0] callResR13;
  logic [130:0] gzdLLziMainzicompute2R6;
  logic [7:0] callResR14;
  logic [130:0] gzdLLziMainzicompute2R7;
  logic [7:0] callResR15;
  logic [63:0] resizzeR9;
  logic [2:0] resizzeR10;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [127:0] resizzeR11;
  logic [2:0] resizzeR12;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [255:0] binOpR14;
  logic [255:0] binOpR15;
  logic [127:0] resizzeR13;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLziMainzicompute7 = {arg0, arg1, arg2, binOpR1[255:128] < binOpR1[127:0]};
  assign gzdLLziMainzicompute6 = {gzdLLziMainzicompute7[131:68], gzdLLziMainzicompute7[67:4], 3'h0};
  zdLLziMainzicompute6  zdLLziMainzicompute6 (gzdLLziMainzicompute6[130:67], gzdLLziMainzicompute6[66:3], gzdLLziMainzicompute6[2:0], callRes);
  assign gzdLLziMainzicompute6R1 = {gzdLLziMainzicompute7[131:68], gzdLLziMainzicompute7[67:4], 3'h1};
  zdLLziMainzicompute6  zdLLziMainzicompute6R1 (gzdLLziMainzicompute6R1[130:67], gzdLLziMainzicompute6R1[66:3], gzdLLziMainzicompute6R1[2:0], callResR1);
  assign gzdLLziMainzicompute6R2 = {gzdLLziMainzicompute7[131:68], gzdLLziMainzicompute7[67:4], 3'h2};
  zdLLziMainzicompute6  zdLLziMainzicompute6R2 (gzdLLziMainzicompute6R2[130:67], gzdLLziMainzicompute6R2[66:3], gzdLLziMainzicompute6R2[2:0], callResR2);
  assign gzdLLziMainzicompute6R3 = {gzdLLziMainzicompute7[131:68], gzdLLziMainzicompute7[67:4], 3'h3};
  zdLLziMainzicompute6  zdLLziMainzicompute6R3 (gzdLLziMainzicompute6R3[130:67], gzdLLziMainzicompute6R3[66:3], gzdLLziMainzicompute6R3[2:0], callResR3);
  assign gzdLLziMainzicompute6R4 = {gzdLLziMainzicompute7[131:68], gzdLLziMainzicompute7[67:4], 3'h4};
  zdLLziMainzicompute6  zdLLziMainzicompute6R4 (gzdLLziMainzicompute6R4[130:67], gzdLLziMainzicompute6R4[66:3], gzdLLziMainzicompute6R4[2:0], callResR4);
  assign gzdLLziMainzicompute6R5 = {gzdLLziMainzicompute7[131:68], gzdLLziMainzicompute7[67:4], 3'h5};
  zdLLziMainzicompute6  zdLLziMainzicompute6R5 (gzdLLziMainzicompute6R5[130:67], gzdLLziMainzicompute6R5[66:3], gzdLLziMainzicompute6R5[2:0], callResR5);
  assign gzdLLziMainzicompute6R6 = {gzdLLziMainzicompute7[131:68], gzdLLziMainzicompute7[67:4], 3'h6};
  zdLLziMainzicompute6  zdLLziMainzicompute6R6 (gzdLLziMainzicompute6R6[130:67], gzdLLziMainzicompute6R6[66:3], gzdLLziMainzicompute6R6[2:0], callResR6);
  assign gzdLLziMainzicompute6R7 = {gzdLLziMainzicompute7[131:68], gzdLLziMainzicompute7[67:4], 3'h7};
  zdLLziMainzicompute6  zdLLziMainzicompute6R7 (gzdLLziMainzicompute6R7[130:67], gzdLLziMainzicompute6R7[66:3], gzdLLziMainzicompute6R7[2:0], callResR7);
  assign resizzeR2 = {callRes, callResR1, callResR2, callResR3, callResR4, callResR5, callResR6, callResR7};
  assign resizzeR3 = gzdLLziMainzicompute7[3:1];
  assign binOpR2 = {128'(resizzeR3[2:0]), 128'h00000000000000000000000000000003};
  assign binOpR3 = {binOpR2[255:128] - binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[2:0];
  assign binOpR4 = {128'(resizzeR5[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR5 = {binOpR4[255:128] * binOpR4[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR6 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR7 = resizzeR6[2:0];
  assign binOpR6 = {128'h00000000000000000000000000000008, 128'(resizzeR7[2:0])};
  assign binOpR7 = {binOpR6[255:128] - binOpR6[127:0], 128'h00000000000000000000000000000001};
  assign binOpR8 = {binOpR7[255:128] - binOpR7[127:0], 128'h00000000000000000000000000000008};
  assign binOpR9 = {128'(resizzeR2[63:0]), binOpR8[255:128] * binOpR8[127:0]};
  assign resizzeR8 = binOpR9[255:128] >> binOpR9[127:0];
  assign gzdLLziMainzicompute3 = {arg0, arg1, arg2, binOp[255:128] < binOp[127:0]};
  assign gzdLLziMainzicompute2 = {gzdLLziMainzicompute3[131:68], gzdLLziMainzicompute3[67:4], 3'h0};
  zdLLziMainzicompute2  zdLLziMainzicompute2 (gzdLLziMainzicompute2[130:67], gzdLLziMainzicompute2[66:3], gzdLLziMainzicompute2[2:0], callResR8);
  assign gzdLLziMainzicompute2R1 = {gzdLLziMainzicompute3[131:68], gzdLLziMainzicompute3[67:4], 3'h1};
  zdLLziMainzicompute2  zdLLziMainzicompute2R1 (gzdLLziMainzicompute2R1[130:67], gzdLLziMainzicompute2R1[66:3], gzdLLziMainzicompute2R1[2:0], callResR9);
  assign gzdLLziMainzicompute2R2 = {gzdLLziMainzicompute3[131:68], gzdLLziMainzicompute3[67:4], 3'h2};
  zdLLziMainzicompute2  zdLLziMainzicompute2R2 (gzdLLziMainzicompute2R2[130:67], gzdLLziMainzicompute2R2[66:3], gzdLLziMainzicompute2R2[2:0], callResR10);
  assign gzdLLziMainzicompute2R3 = {gzdLLziMainzicompute3[131:68], gzdLLziMainzicompute3[67:4], 3'h3};
  zdLLziMainzicompute2  zdLLziMainzicompute2R3 (gzdLLziMainzicompute2R3[130:67], gzdLLziMainzicompute2R3[66:3], gzdLLziMainzicompute2R3[2:0], callResR11);
  assign gzdLLziMainzicompute2R4 = {gzdLLziMainzicompute3[131:68], gzdLLziMainzicompute3[67:4], 3'h4};
  zdLLziMainzicompute2  zdLLziMainzicompute2R4 (gzdLLziMainzicompute2R4[130:67], gzdLLziMainzicompute2R4[66:3], gzdLLziMainzicompute2R4[2:0], callResR12);
  assign gzdLLziMainzicompute2R5 = {gzdLLziMainzicompute3[131:68], gzdLLziMainzicompute3[67:4], 3'h5};
  zdLLziMainzicompute2  zdLLziMainzicompute2R5 (gzdLLziMainzicompute2R5[130:67], gzdLLziMainzicompute2R5[66:3], gzdLLziMainzicompute2R5[2:0], callResR13);
  assign gzdLLziMainzicompute2R6 = {gzdLLziMainzicompute3[131:68], gzdLLziMainzicompute3[67:4], 3'h6};
  zdLLziMainzicompute2  zdLLziMainzicompute2R6 (gzdLLziMainzicompute2R6[130:67], gzdLLziMainzicompute2R6[66:3], gzdLLziMainzicompute2R6[2:0], callResR14);
  assign gzdLLziMainzicompute2R7 = {gzdLLziMainzicompute3[131:68], gzdLLziMainzicompute3[67:4], 3'h7};
  zdLLziMainzicompute2  zdLLziMainzicompute2R7 (gzdLLziMainzicompute2R7[130:67], gzdLLziMainzicompute2R7[66:3], gzdLLziMainzicompute2R7[2:0], callResR15);
  assign resizzeR9 = {callResR8, callResR9, callResR10, callResR11, callResR12, callResR13, callResR14, callResR15};
  assign resizzeR10 = gzdLLziMainzicompute3[3:1];
  assign binOpR10 = {128'(resizzeR10[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR11 = {binOpR10[255:128] * binOpR10[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR11 = binOpR11[255:128] % binOpR11[127:0];
  assign resizzeR12 = resizzeR11[2:0];
  assign binOpR12 = {128'h00000000000000000000000000000008, 128'(resizzeR12[2:0])};
  assign binOpR13 = {binOpR12[255:128] - binOpR12[127:0], 128'h00000000000000000000000000000001};
  assign binOpR14 = {binOpR13[255:128] - binOpR13[127:0], 128'h00000000000000000000000000000008};
  assign binOpR15 = {128'(resizzeR9[63:0]), binOpR14[255:128] * binOpR14[127:0]};
  assign resizzeR13 = binOpR15[255:128] >> binOpR15[127:0];
  assign res = (gzdLLziMainzicompute3[0] == 1'h1) ? resizzeR13[7:0] : resizzeR8[7:0];
endmodule

module zdLLziMainzicompute12 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [67:0] gzdLLziMainzicompute1;
  logic [7:0] callRes;
  logic [67:0] gzdLLziMainzicompute;
  logic [7:0] callResR1;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLziMainzicompute1 = {arg1, arg2, binOpR1[255:128] < binOpR1[127:0]};
  zdLLziMainzicompute1  zdLLziMainzicompute1 (gzdLLziMainzicompute1[67:4], gzdLLziMainzicompute1[3:1], callRes);
  assign gzdLLziMainzicompute = {arg0, arg2, binOp[255:128] < binOp[127:0]};
  zdLLziMainzicompute  zdLLziMainzicompute (gzdLLziMainzicompute[67:4], gzdLLziMainzicompute[3:1], callResR1);
  assign res = (gzdLLziMainzicompute[0] == 1'h1) ? callResR1 : callRes;
endmodule

module zdLLziMainzicompute14 (input logic [63:0] arg0,
  input logic [2:0] arg1,
  output logic [7:0] res);
  logic [63:0] resizze;
  logic [2:0] resizzeR1;
  logic [255:0] binOp;
  logic [255:0] binOpR1;
  logic [127:0] resizzeR2;
  logic [2:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR4;
  assign resizze = arg0;
  assign resizzeR1 = arg1;
  assign binOp = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR1 = {binOp[255:128] * binOp[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR2 = binOpR1[255:128] % binOpR1[127:0];
  assign resizzeR3 = resizzeR2[2:0];
  assign binOpR2 = {128'h00000000000000000000000000000008, 128'(resizzeR3[2:0])};
  assign binOpR3 = {binOpR2[255:128] - binOpR2[127:0], 128'h00000000000000000000000000000001};
  assign binOpR4 = {binOpR3[255:128] - binOpR3[127:0], 128'h00000000000000000000000000000008};
  assign binOpR5 = {128'(resizze[63:0]), binOpR4[255:128] * binOpR4[127:0]};
  assign resizzeR4 = binOpR5[255:128] >> binOpR5[127:0];
  assign res = resizzeR4[7:0];
endmodule

module zdLLziMainzicompute15 (input logic [63:0] arg0,
  input logic [2:0] arg1,
  output logic [7:0] res);
  logic [63:0] resizze;
  logic [2:0] resizzeR1;
  logic [255:0] binOp;
  logic [255:0] binOpR1;
  logic [127:0] resizzeR2;
  logic [2:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [127:0] resizzeR6;
  assign resizze = arg0;
  assign resizzeR1 = arg1;
  assign binOp = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign binOpR1 = {binOp[255:128] - binOp[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR2 = binOpR1[255:128] % binOpR1[127:0];
  assign resizzeR3 = resizzeR2[2:0];
  assign binOpR2 = {128'(resizzeR3[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR3 = {binOpR2[255:128] * binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[2:0];
  assign binOpR4 = {128'h00000000000000000000000000000008, 128'(resizzeR5[2:0])};
  assign binOpR5 = {binOpR4[255:128] - binOpR4[127:0], 128'h00000000000000000000000000000001};
  assign binOpR6 = {binOpR5[255:128] - binOpR5[127:0], 128'h00000000000000000000000000000008};
  assign binOpR7 = {128'(resizze[63:0]), binOpR6[255:128] * binOpR6[127:0]};
  assign resizzeR6 = binOpR7[255:128] >> binOpR7[127:0];
  assign res = resizzeR6[7:0];
endmodule

module zdLLziMainzicompute16 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [67:0] gzdLLziMainzicompute15;
  logic [7:0] callRes;
  logic [67:0] gzdLLziMainzicompute14;
  logic [7:0] callResR1;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLziMainzicompute15 = {arg1, arg2, binOpR1[255:128] < binOpR1[127:0]};
  zdLLziMainzicompute15  zdLLziMainzicompute15 (gzdLLziMainzicompute15[67:4], gzdLLziMainzicompute15[3:1], callRes);
  assign gzdLLziMainzicompute14 = {arg0, arg2, binOp[255:128] < binOp[127:0]};
  zdLLziMainzicompute14  zdLLziMainzicompute14 (gzdLLziMainzicompute14[67:4], gzdLLziMainzicompute14[3:1], callResR1);
  assign res = (gzdLLziMainzicompute14[0] == 1'h1) ? callResR1 : callRes;
endmodule

module zdLLziMainzicompute18 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [131:0] gzdLLziMainzicompute17;
  logic [130:0] gzdLLziMainzicompute16;
  logic [7:0] callRes;
  logic [130:0] gzdLLziMainzicompute16R1;
  logic [7:0] callResR1;
  logic [130:0] gzdLLziMainzicompute16R2;
  logic [7:0] callResR2;
  logic [130:0] gzdLLziMainzicompute16R3;
  logic [7:0] callResR3;
  logic [130:0] gzdLLziMainzicompute16R4;
  logic [7:0] callResR4;
  logic [130:0] gzdLLziMainzicompute16R5;
  logic [7:0] callResR5;
  logic [130:0] gzdLLziMainzicompute16R6;
  logic [7:0] callResR6;
  logic [130:0] gzdLLziMainzicompute16R7;
  logic [7:0] callResR7;
  logic [63:0] resizzeR2;
  logic [2:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR6;
  logic [2:0] resizzeR7;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [127:0] resizzeR8;
  logic [2:0] resizzeR9;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [127:0] resizzeR10;
  logic [131:0] gzdLLziMainzicompute13;
  logic [130:0] gzdLLziMainzicompute12;
  logic [7:0] callResR8;
  logic [130:0] gzdLLziMainzicompute12R1;
  logic [7:0] callResR9;
  logic [130:0] gzdLLziMainzicompute12R2;
  logic [7:0] callResR10;
  logic [130:0] gzdLLziMainzicompute12R3;
  logic [7:0] callResR11;
  logic [130:0] gzdLLziMainzicompute12R4;
  logic [7:0] callResR12;
  logic [130:0] gzdLLziMainzicompute12R5;
  logic [7:0] callResR13;
  logic [130:0] gzdLLziMainzicompute12R6;
  logic [7:0] callResR14;
  logic [130:0] gzdLLziMainzicompute12R7;
  logic [7:0] callResR15;
  logic [63:0] resizzeR11;
  logic [2:0] resizzeR12;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [127:0] resizzeR13;
  logic [2:0] resizzeR14;
  logic [255:0] binOpR14;
  logic [255:0] binOpR15;
  logic [127:0] resizzeR15;
  logic [2:0] resizzeR16;
  logic [255:0] binOpR16;
  logic [255:0] binOpR17;
  logic [255:0] binOpR18;
  logic [255:0] binOpR19;
  logic [127:0] resizzeR17;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLziMainzicompute17 = {arg0, arg1, arg2, binOpR1[255:128] < binOpR1[127:0]};
  assign gzdLLziMainzicompute16 = {gzdLLziMainzicompute17[131:68], gzdLLziMainzicompute17[67:4], 3'h0};
  zdLLziMainzicompute16  zdLLziMainzicompute16 (gzdLLziMainzicompute16[130:67], gzdLLziMainzicompute16[66:3], gzdLLziMainzicompute16[2:0], callRes);
  assign gzdLLziMainzicompute16R1 = {gzdLLziMainzicompute17[131:68], gzdLLziMainzicompute17[67:4], 3'h1};
  zdLLziMainzicompute16  zdLLziMainzicompute16R1 (gzdLLziMainzicompute16R1[130:67], gzdLLziMainzicompute16R1[66:3], gzdLLziMainzicompute16R1[2:0], callResR1);
  assign gzdLLziMainzicompute16R2 = {gzdLLziMainzicompute17[131:68], gzdLLziMainzicompute17[67:4], 3'h2};
  zdLLziMainzicompute16  zdLLziMainzicompute16R2 (gzdLLziMainzicompute16R2[130:67], gzdLLziMainzicompute16R2[66:3], gzdLLziMainzicompute16R2[2:0], callResR2);
  assign gzdLLziMainzicompute16R3 = {gzdLLziMainzicompute17[131:68], gzdLLziMainzicompute17[67:4], 3'h3};
  zdLLziMainzicompute16  zdLLziMainzicompute16R3 (gzdLLziMainzicompute16R3[130:67], gzdLLziMainzicompute16R3[66:3], gzdLLziMainzicompute16R3[2:0], callResR3);
  assign gzdLLziMainzicompute16R4 = {gzdLLziMainzicompute17[131:68], gzdLLziMainzicompute17[67:4], 3'h4};
  zdLLziMainzicompute16  zdLLziMainzicompute16R4 (gzdLLziMainzicompute16R4[130:67], gzdLLziMainzicompute16R4[66:3], gzdLLziMainzicompute16R4[2:0], callResR4);
  assign gzdLLziMainzicompute16R5 = {gzdLLziMainzicompute17[131:68], gzdLLziMainzicompute17[67:4], 3'h5};
  zdLLziMainzicompute16  zdLLziMainzicompute16R5 (gzdLLziMainzicompute16R5[130:67], gzdLLziMainzicompute16R5[66:3], gzdLLziMainzicompute16R5[2:0], callResR5);
  assign gzdLLziMainzicompute16R6 = {gzdLLziMainzicompute17[131:68], gzdLLziMainzicompute17[67:4], 3'h6};
  zdLLziMainzicompute16  zdLLziMainzicompute16R6 (gzdLLziMainzicompute16R6[130:67], gzdLLziMainzicompute16R6[66:3], gzdLLziMainzicompute16R6[2:0], callResR6);
  assign gzdLLziMainzicompute16R7 = {gzdLLziMainzicompute17[131:68], gzdLLziMainzicompute17[67:4], 3'h7};
  zdLLziMainzicompute16  zdLLziMainzicompute16R7 (gzdLLziMainzicompute16R7[130:67], gzdLLziMainzicompute16R7[66:3], gzdLLziMainzicompute16R7[2:0], callResR7);
  assign resizzeR2 = {callRes, callResR1, callResR2, callResR3, callResR4, callResR5, callResR6, callResR7};
  assign resizzeR3 = gzdLLziMainzicompute17[3:1];
  assign binOpR2 = {128'(resizzeR3[2:0]), 128'h00000000000000000000000000000003};
  assign binOpR3 = {binOpR2[255:128] - binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[2:0];
  assign binOpR4 = {128'(resizzeR5[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR5 = {binOpR4[255:128] * binOpR4[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR6 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR7 = resizzeR6[2:0];
  assign binOpR6 = {128'(resizzeR7[2:0]), 128'h00000000000000000000000000000001};
  assign binOpR7 = {binOpR6[255:128] + binOpR6[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR8 = binOpR7[255:128] % binOpR7[127:0];
  assign resizzeR9 = resizzeR8[2:0];
  assign binOpR8 = {128'h00000000000000000000000000000008, 128'(resizzeR9[2:0])};
  assign binOpR9 = {binOpR8[255:128] - binOpR8[127:0], 128'h00000000000000000000000000000001};
  assign binOpR10 = {binOpR9[255:128] - binOpR9[127:0], 128'h00000000000000000000000000000008};
  assign binOpR11 = {128'(resizzeR2[63:0]), binOpR10[255:128] * binOpR10[127:0]};
  assign resizzeR10 = binOpR11[255:128] >> binOpR11[127:0];
  assign gzdLLziMainzicompute13 = {arg0, arg1, arg2, binOp[255:128] < binOp[127:0]};
  assign gzdLLziMainzicompute12 = {gzdLLziMainzicompute13[131:68], gzdLLziMainzicompute13[67:4], 3'h0};
  zdLLziMainzicompute12  zdLLziMainzicompute12 (gzdLLziMainzicompute12[130:67], gzdLLziMainzicompute12[66:3], gzdLLziMainzicompute12[2:0], callResR8);
  assign gzdLLziMainzicompute12R1 = {gzdLLziMainzicompute13[131:68], gzdLLziMainzicompute13[67:4], 3'h1};
  zdLLziMainzicompute12  zdLLziMainzicompute12R1 (gzdLLziMainzicompute12R1[130:67], gzdLLziMainzicompute12R1[66:3], gzdLLziMainzicompute12R1[2:0], callResR9);
  assign gzdLLziMainzicompute12R2 = {gzdLLziMainzicompute13[131:68], gzdLLziMainzicompute13[67:4], 3'h2};
  zdLLziMainzicompute12  zdLLziMainzicompute12R2 (gzdLLziMainzicompute12R2[130:67], gzdLLziMainzicompute12R2[66:3], gzdLLziMainzicompute12R2[2:0], callResR10);
  assign gzdLLziMainzicompute12R3 = {gzdLLziMainzicompute13[131:68], gzdLLziMainzicompute13[67:4], 3'h3};
  zdLLziMainzicompute12  zdLLziMainzicompute12R3 (gzdLLziMainzicompute12R3[130:67], gzdLLziMainzicompute12R3[66:3], gzdLLziMainzicompute12R3[2:0], callResR11);
  assign gzdLLziMainzicompute12R4 = {gzdLLziMainzicompute13[131:68], gzdLLziMainzicompute13[67:4], 3'h4};
  zdLLziMainzicompute12  zdLLziMainzicompute12R4 (gzdLLziMainzicompute12R4[130:67], gzdLLziMainzicompute12R4[66:3], gzdLLziMainzicompute12R4[2:0], callResR12);
  assign gzdLLziMainzicompute12R5 = {gzdLLziMainzicompute13[131:68], gzdLLziMainzicompute13[67:4], 3'h5};
  zdLLziMainzicompute12  zdLLziMainzicompute12R5 (gzdLLziMainzicompute12R5[130:67], gzdLLziMainzicompute12R5[66:3], gzdLLziMainzicompute12R5[2:0], callResR13);
  assign gzdLLziMainzicompute12R6 = {gzdLLziMainzicompute13[131:68], gzdLLziMainzicompute13[67:4], 3'h6};
  zdLLziMainzicompute12  zdLLziMainzicompute12R6 (gzdLLziMainzicompute12R6[130:67], gzdLLziMainzicompute12R6[66:3], gzdLLziMainzicompute12R6[2:0], callResR14);
  assign gzdLLziMainzicompute12R7 = {gzdLLziMainzicompute13[131:68], gzdLLziMainzicompute13[67:4], 3'h7};
  zdLLziMainzicompute12  zdLLziMainzicompute12R7 (gzdLLziMainzicompute12R7[130:67], gzdLLziMainzicompute12R7[66:3], gzdLLziMainzicompute12R7[2:0], callResR15);
  assign resizzeR11 = {callResR8, callResR9, callResR10, callResR11, callResR12, callResR13, callResR14, callResR15};
  assign resizzeR12 = gzdLLziMainzicompute13[3:1];
  assign binOpR12 = {128'(resizzeR12[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR13 = {binOpR12[255:128] * binOpR12[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR13 = binOpR13[255:128] % binOpR13[127:0];
  assign resizzeR14 = resizzeR13[2:0];
  assign binOpR14 = {128'(resizzeR14[2:0]), 128'h00000000000000000000000000000001};
  assign binOpR15 = {binOpR14[255:128] + binOpR14[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR15 = binOpR15[255:128] % binOpR15[127:0];
  assign resizzeR16 = resizzeR15[2:0];
  assign binOpR16 = {128'h00000000000000000000000000000008, 128'(resizzeR16[2:0])};
  assign binOpR17 = {binOpR16[255:128] - binOpR16[127:0], 128'h00000000000000000000000000000001};
  assign binOpR18 = {binOpR17[255:128] - binOpR17[127:0], 128'h00000000000000000000000000000008};
  assign binOpR19 = {128'(resizzeR11[63:0]), binOpR18[255:128] * binOpR18[127:0]};
  assign resizzeR17 = binOpR19[255:128] >> binOpR19[127:0];
  assign res = (gzdLLziMainzicompute13[0] == 1'h1) ? resizzeR17[7:0] : resizzeR10[7:0];
endmodule

module zdLLziMainzicompute20 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [127:0] resizzeR1;
  logic [0:0] msbit;
  logic [0:0] gReWireziPreludezinot;
  logic [0:0] callRes;
  logic [2:0] resizzeR2;
  logic [127:0] resizzeR3;
  logic [0:0] msbitR1;
  logic [0:0] gReWireziPreludezinotR1;
  logic [0:0] callResR1;
  logic [131:0] gzdLLziMainzicompute19;
  logic [130:0] gzdLLziMainzicompute18;
  logic [7:0] callResR2;
  logic [130:0] gzdLLziMainzicompute18R1;
  logic [7:0] callResR3;
  logic [130:0] gzdLLziMainzicompute18R2;
  logic [7:0] callResR4;
  logic [130:0] gzdLLziMainzicompute18R3;
  logic [7:0] callResR5;
  logic [130:0] gzdLLziMainzicompute18R4;
  logic [7:0] callResR6;
  logic [130:0] gzdLLziMainzicompute18R5;
  logic [7:0] callResR7;
  logic [130:0] gzdLLziMainzicompute18R6;
  logic [7:0] callResR8;
  logic [130:0] gzdLLziMainzicompute18R7;
  logic [7:0] callResR9;
  logic [63:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOp;
  logic [255:0] binOpR1;
  logic [127:0] resizzeR6;
  logic [2:0] resizzeR7;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR8;
  logic [2:0] resizzeR9;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [127:0] resizzeR10;
  logic [131:0] gzdLLziMainzicompute9;
  logic [130:0] gzdLLziMainzicompute8;
  logic [7:0] callResR10;
  logic [130:0] gzdLLziMainzicompute8R1;
  logic [7:0] callResR11;
  logic [130:0] gzdLLziMainzicompute8R2;
  logic [7:0] callResR12;
  logic [130:0] gzdLLziMainzicompute8R3;
  logic [7:0] callResR13;
  logic [130:0] gzdLLziMainzicompute8R4;
  logic [7:0] callResR14;
  logic [130:0] gzdLLziMainzicompute8R5;
  logic [7:0] callResR15;
  logic [130:0] gzdLLziMainzicompute8R6;
  logic [7:0] callResR16;
  logic [130:0] gzdLLziMainzicompute8R7;
  logic [7:0] callResR17;
  logic [63:0] resizzeR11;
  logic [2:0] resizzeR12;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [127:0] resizzeR13;
  logic [2:0] resizzeR14;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [127:0] resizzeR15;
  assign resizze = arg2;
  assign resizzeR1 = 128'(resizze[2:0]);
  assign msbit = resizzeR1[0];
  assign gReWireziPreludezinot = msbit[0];
  ReWireziPreludezinot  ReWireziPreludezinot (gReWireziPreludezinot[0], callRes);
  assign resizzeR2 = arg2;
  assign resizzeR3 = 128'(resizzeR2[2:0]);
  assign msbitR1 = resizzeR3[0];
  assign gReWireziPreludezinotR1 = msbitR1[0];
  ReWireziPreludezinot  ReWireziPreludezinotR1 (gReWireziPreludezinotR1[0], callResR1);
  assign gzdLLziMainzicompute19 = {arg0, arg1, arg2, callResR1};
  assign gzdLLziMainzicompute18 = {gzdLLziMainzicompute19[131:68], gzdLLziMainzicompute19[67:4], 3'h0};
  zdLLziMainzicompute18  zdLLziMainzicompute18 (gzdLLziMainzicompute18[130:67], gzdLLziMainzicompute18[66:3], gzdLLziMainzicompute18[2:0], callResR2);
  assign gzdLLziMainzicompute18R1 = {gzdLLziMainzicompute19[131:68], gzdLLziMainzicompute19[67:4], 3'h1};
  zdLLziMainzicompute18  zdLLziMainzicompute18R1 (gzdLLziMainzicompute18R1[130:67], gzdLLziMainzicompute18R1[66:3], gzdLLziMainzicompute18R1[2:0], callResR3);
  assign gzdLLziMainzicompute18R2 = {gzdLLziMainzicompute19[131:68], gzdLLziMainzicompute19[67:4], 3'h2};
  zdLLziMainzicompute18  zdLLziMainzicompute18R2 (gzdLLziMainzicompute18R2[130:67], gzdLLziMainzicompute18R2[66:3], gzdLLziMainzicompute18R2[2:0], callResR4);
  assign gzdLLziMainzicompute18R3 = {gzdLLziMainzicompute19[131:68], gzdLLziMainzicompute19[67:4], 3'h3};
  zdLLziMainzicompute18  zdLLziMainzicompute18R3 (gzdLLziMainzicompute18R3[130:67], gzdLLziMainzicompute18R3[66:3], gzdLLziMainzicompute18R3[2:0], callResR5);
  assign gzdLLziMainzicompute18R4 = {gzdLLziMainzicompute19[131:68], gzdLLziMainzicompute19[67:4], 3'h4};
  zdLLziMainzicompute18  zdLLziMainzicompute18R4 (gzdLLziMainzicompute18R4[130:67], gzdLLziMainzicompute18R4[66:3], gzdLLziMainzicompute18R4[2:0], callResR6);
  assign gzdLLziMainzicompute18R5 = {gzdLLziMainzicompute19[131:68], gzdLLziMainzicompute19[67:4], 3'h5};
  zdLLziMainzicompute18  zdLLziMainzicompute18R5 (gzdLLziMainzicompute18R5[130:67], gzdLLziMainzicompute18R5[66:3], gzdLLziMainzicompute18R5[2:0], callResR7);
  assign gzdLLziMainzicompute18R6 = {gzdLLziMainzicompute19[131:68], gzdLLziMainzicompute19[67:4], 3'h6};
  zdLLziMainzicompute18  zdLLziMainzicompute18R6 (gzdLLziMainzicompute18R6[130:67], gzdLLziMainzicompute18R6[66:3], gzdLLziMainzicompute18R6[2:0], callResR8);
  assign gzdLLziMainzicompute18R7 = {gzdLLziMainzicompute19[131:68], gzdLLziMainzicompute19[67:4], 3'h7};
  zdLLziMainzicompute18  zdLLziMainzicompute18R7 (gzdLLziMainzicompute18R7[130:67], gzdLLziMainzicompute18R7[66:3], gzdLLziMainzicompute18R7[2:0], callResR9);
  assign resizzeR4 = {callResR2, callResR3, callResR4, callResR5, callResR6, callResR7, callResR8, callResR9};
  assign resizzeR5 = gzdLLziMainzicompute19[3:1];
  assign binOp = {128'(resizzeR5[2:0]), 128'h00000000000000000000000000000001};
  assign binOpR1 = {binOp[255:128] - binOp[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR6 = binOpR1[255:128] % binOpR1[127:0];
  assign resizzeR7 = resizzeR6[2:0];
  assign binOpR2 = {128'(resizzeR7[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR3 = {binOpR2[255:128] / binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR8 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR9 = resizzeR8[2:0];
  assign binOpR4 = {128'h00000000000000000000000000000008, 128'(resizzeR9[2:0])};
  assign binOpR5 = {binOpR4[255:128] - binOpR4[127:0], 128'h00000000000000000000000000000001};
  assign binOpR6 = {binOpR5[255:128] - binOpR5[127:0], 128'h00000000000000000000000000000008};
  assign binOpR7 = {128'(resizzeR4[63:0]), binOpR6[255:128] * binOpR6[127:0]};
  assign resizzeR10 = binOpR7[255:128] >> binOpR7[127:0];
  assign gzdLLziMainzicompute9 = {arg0, arg1, arg2, callRes};
  assign gzdLLziMainzicompute8 = {gzdLLziMainzicompute9[131:68], gzdLLziMainzicompute9[67:4], 3'h0};
  zdLLziMainzicompute8  zdLLziMainzicompute8 (gzdLLziMainzicompute8[130:67], gzdLLziMainzicompute8[66:3], gzdLLziMainzicompute8[2:0], callResR10);
  assign gzdLLziMainzicompute8R1 = {gzdLLziMainzicompute9[131:68], gzdLLziMainzicompute9[67:4], 3'h1};
  zdLLziMainzicompute8  zdLLziMainzicompute8R1 (gzdLLziMainzicompute8R1[130:67], gzdLLziMainzicompute8R1[66:3], gzdLLziMainzicompute8R1[2:0], callResR11);
  assign gzdLLziMainzicompute8R2 = {gzdLLziMainzicompute9[131:68], gzdLLziMainzicompute9[67:4], 3'h2};
  zdLLziMainzicompute8  zdLLziMainzicompute8R2 (gzdLLziMainzicompute8R2[130:67], gzdLLziMainzicompute8R2[66:3], gzdLLziMainzicompute8R2[2:0], callResR12);
  assign gzdLLziMainzicompute8R3 = {gzdLLziMainzicompute9[131:68], gzdLLziMainzicompute9[67:4], 3'h3};
  zdLLziMainzicompute8  zdLLziMainzicompute8R3 (gzdLLziMainzicompute8R3[130:67], gzdLLziMainzicompute8R3[66:3], gzdLLziMainzicompute8R3[2:0], callResR13);
  assign gzdLLziMainzicompute8R4 = {gzdLLziMainzicompute9[131:68], gzdLLziMainzicompute9[67:4], 3'h4};
  zdLLziMainzicompute8  zdLLziMainzicompute8R4 (gzdLLziMainzicompute8R4[130:67], gzdLLziMainzicompute8R4[66:3], gzdLLziMainzicompute8R4[2:0], callResR14);
  assign gzdLLziMainzicompute8R5 = {gzdLLziMainzicompute9[131:68], gzdLLziMainzicompute9[67:4], 3'h5};
  zdLLziMainzicompute8  zdLLziMainzicompute8R5 (gzdLLziMainzicompute8R5[130:67], gzdLLziMainzicompute8R5[66:3], gzdLLziMainzicompute8R5[2:0], callResR15);
  assign gzdLLziMainzicompute8R6 = {gzdLLziMainzicompute9[131:68], gzdLLziMainzicompute9[67:4], 3'h6};
  zdLLziMainzicompute8  zdLLziMainzicompute8R6 (gzdLLziMainzicompute8R6[130:67], gzdLLziMainzicompute8R6[66:3], gzdLLziMainzicompute8R6[2:0], callResR16);
  assign gzdLLziMainzicompute8R7 = {gzdLLziMainzicompute9[131:68], gzdLLziMainzicompute9[67:4], 3'h7};
  zdLLziMainzicompute8  zdLLziMainzicompute8R7 (gzdLLziMainzicompute8R7[130:67], gzdLLziMainzicompute8R7[66:3], gzdLLziMainzicompute8R7[2:0], callResR17);
  assign resizzeR11 = {callResR10, callResR11, callResR12, callResR13, callResR14, callResR15, callResR16, callResR17};
  assign resizzeR12 = gzdLLziMainzicompute9[3:1];
  assign binOpR8 = {128'(resizzeR12[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR9 = {binOpR8[255:128] / binOpR8[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR13 = binOpR9[255:128] % binOpR9[127:0];
  assign resizzeR14 = resizzeR13[2:0];
  assign binOpR10 = {128'h00000000000000000000000000000008, 128'(resizzeR14[2:0])};
  assign binOpR11 = {binOpR10[255:128] - binOpR10[127:0], 128'h00000000000000000000000000000001};
  assign binOpR12 = {binOpR11[255:128] - binOpR11[127:0], 128'h00000000000000000000000000000008};
  assign binOpR13 = {128'(resizzeR11[63:0]), binOpR12[255:128] * binOpR12[127:0]};
  assign resizzeR15 = binOpR13[255:128] >> binOpR13[127:0];
  assign res = (gzdLLziMainzicompute9[0] == 1'h1) ? resizzeR15[7:0] : resizzeR10[7:0];
endmodule

module zdLLziMainzicompute23 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [67:0] gzdLLziMainzicompute1;
  logic [7:0] callRes;
  logic [67:0] gzdLLziMainzicompute;
  logic [7:0] callResR1;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLziMainzicompute1 = {arg1, arg2, binOpR1[255:128] < binOpR1[127:0]};
  zdLLziMainzicompute1  zdLLziMainzicompute1 (gzdLLziMainzicompute1[67:4], gzdLLziMainzicompute1[3:1], callRes);
  assign gzdLLziMainzicompute = {arg0, arg2, binOp[255:128] < binOp[127:0]};
  zdLLziMainzicompute  zdLLziMainzicompute (gzdLLziMainzicompute[67:4], gzdLLziMainzicompute[3:1], callResR1);
  assign res = (gzdLLziMainzicompute[0] == 1'h1) ? callResR1 : callRes;
endmodule

module zdLLziMainzicompute27 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [67:0] gzdLLziMainzicompute15;
  logic [7:0] callRes;
  logic [67:0] gzdLLziMainzicompute14;
  logic [7:0] callResR1;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLziMainzicompute15 = {arg1, arg2, binOpR1[255:128] < binOpR1[127:0]};
  zdLLziMainzicompute15  zdLLziMainzicompute15 (gzdLLziMainzicompute15[67:4], gzdLLziMainzicompute15[3:1], callRes);
  assign gzdLLziMainzicompute14 = {arg0, arg2, binOp[255:128] < binOp[127:0]};
  zdLLziMainzicompute14  zdLLziMainzicompute14 (gzdLLziMainzicompute14[67:4], gzdLLziMainzicompute14[3:1], callResR1);
  assign res = (gzdLLziMainzicompute14[0] == 1'h1) ? callResR1 : callRes;
endmodule

module zdLLziMainzicompute29 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [131:0] gzdLLziMainzicompute28;
  logic [130:0] gzdLLziMainzicompute27;
  logic [7:0] callRes;
  logic [130:0] gzdLLziMainzicompute27R1;
  logic [7:0] callResR1;
  logic [130:0] gzdLLziMainzicompute27R2;
  logic [7:0] callResR2;
  logic [130:0] gzdLLziMainzicompute27R3;
  logic [7:0] callResR3;
  logic [130:0] gzdLLziMainzicompute27R4;
  logic [7:0] callResR4;
  logic [130:0] gzdLLziMainzicompute27R5;
  logic [7:0] callResR5;
  logic [130:0] gzdLLziMainzicompute27R6;
  logic [7:0] callResR6;
  logic [130:0] gzdLLziMainzicompute27R7;
  logic [7:0] callResR7;
  logic [63:0] resizzeR2;
  logic [2:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR6;
  logic [2:0] resizzeR7;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [127:0] resizzeR8;
  logic [131:0] gzdLLziMainzicompute24;
  logic [130:0] gzdLLziMainzicompute23;
  logic [7:0] callResR8;
  logic [130:0] gzdLLziMainzicompute23R1;
  logic [7:0] callResR9;
  logic [130:0] gzdLLziMainzicompute23R2;
  logic [7:0] callResR10;
  logic [130:0] gzdLLziMainzicompute23R3;
  logic [7:0] callResR11;
  logic [130:0] gzdLLziMainzicompute23R4;
  logic [7:0] callResR12;
  logic [130:0] gzdLLziMainzicompute23R5;
  logic [7:0] callResR13;
  logic [130:0] gzdLLziMainzicompute23R6;
  logic [7:0] callResR14;
  logic [130:0] gzdLLziMainzicompute23R7;
  logic [7:0] callResR15;
  logic [63:0] resizzeR9;
  logic [2:0] resizzeR10;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [127:0] resizzeR11;
  logic [2:0] resizzeR12;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [255:0] binOpR14;
  logic [255:0] binOpR15;
  logic [127:0] resizzeR13;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLziMainzicompute28 = {arg2, arg0, arg1, binOpR1[255:128] < binOpR1[127:0]};
  assign gzdLLziMainzicompute27 = {gzdLLziMainzicompute28[128:65], gzdLLziMainzicompute28[64:1], 3'h0};
  zdLLziMainzicompute27  zdLLziMainzicompute27 (gzdLLziMainzicompute27[130:67], gzdLLziMainzicompute27[66:3], gzdLLziMainzicompute27[2:0], callRes);
  assign gzdLLziMainzicompute27R1 = {gzdLLziMainzicompute28[128:65], gzdLLziMainzicompute28[64:1], 3'h1};
  zdLLziMainzicompute27  zdLLziMainzicompute27R1 (gzdLLziMainzicompute27R1[130:67], gzdLLziMainzicompute27R1[66:3], gzdLLziMainzicompute27R1[2:0], callResR1);
  assign gzdLLziMainzicompute27R2 = {gzdLLziMainzicompute28[128:65], gzdLLziMainzicompute28[64:1], 3'h2};
  zdLLziMainzicompute27  zdLLziMainzicompute27R2 (gzdLLziMainzicompute27R2[130:67], gzdLLziMainzicompute27R2[66:3], gzdLLziMainzicompute27R2[2:0], callResR2);
  assign gzdLLziMainzicompute27R3 = {gzdLLziMainzicompute28[128:65], gzdLLziMainzicompute28[64:1], 3'h3};
  zdLLziMainzicompute27  zdLLziMainzicompute27R3 (gzdLLziMainzicompute27R3[130:67], gzdLLziMainzicompute27R3[66:3], gzdLLziMainzicompute27R3[2:0], callResR3);
  assign gzdLLziMainzicompute27R4 = {gzdLLziMainzicompute28[128:65], gzdLLziMainzicompute28[64:1], 3'h4};
  zdLLziMainzicompute27  zdLLziMainzicompute27R4 (gzdLLziMainzicompute27R4[130:67], gzdLLziMainzicompute27R4[66:3], gzdLLziMainzicompute27R4[2:0], callResR4);
  assign gzdLLziMainzicompute27R5 = {gzdLLziMainzicompute28[128:65], gzdLLziMainzicompute28[64:1], 3'h5};
  zdLLziMainzicompute27  zdLLziMainzicompute27R5 (gzdLLziMainzicompute27R5[130:67], gzdLLziMainzicompute27R5[66:3], gzdLLziMainzicompute27R5[2:0], callResR5);
  assign gzdLLziMainzicompute27R6 = {gzdLLziMainzicompute28[128:65], gzdLLziMainzicompute28[64:1], 3'h6};
  zdLLziMainzicompute27  zdLLziMainzicompute27R6 (gzdLLziMainzicompute27R6[130:67], gzdLLziMainzicompute27R6[66:3], gzdLLziMainzicompute27R6[2:0], callResR6);
  assign gzdLLziMainzicompute27R7 = {gzdLLziMainzicompute28[128:65], gzdLLziMainzicompute28[64:1], 3'h7};
  zdLLziMainzicompute27  zdLLziMainzicompute27R7 (gzdLLziMainzicompute27R7[130:67], gzdLLziMainzicompute27R7[66:3], gzdLLziMainzicompute27R7[2:0], callResR7);
  assign resizzeR2 = {callRes, callResR1, callResR2, callResR3, callResR4, callResR5, callResR6, callResR7};
  assign resizzeR3 = gzdLLziMainzicompute28[131:129];
  assign binOpR2 = {128'(resizzeR3[2:0]), 128'h00000000000000000000000000000003};
  assign binOpR3 = {binOpR2[255:128] - binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[2:0];
  assign binOpR4 = {128'(resizzeR5[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR5 = {binOpR4[255:128] * binOpR4[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR6 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR7 = resizzeR6[2:0];
  assign binOpR6 = {128'h00000000000000000000000000000008, 128'(resizzeR7[2:0])};
  assign binOpR7 = {binOpR6[255:128] - binOpR6[127:0], 128'h00000000000000000000000000000001};
  assign binOpR8 = {binOpR7[255:128] - binOpR7[127:0], 128'h00000000000000000000000000000008};
  assign binOpR9 = {128'(resizzeR2[63:0]), binOpR8[255:128] * binOpR8[127:0]};
  assign resizzeR8 = binOpR9[255:128] >> binOpR9[127:0];
  assign gzdLLziMainzicompute24 = {arg2, arg0, arg1, binOp[255:128] < binOp[127:0]};
  assign gzdLLziMainzicompute23 = {gzdLLziMainzicompute24[128:65], gzdLLziMainzicompute24[64:1], 3'h0};
  zdLLziMainzicompute23  zdLLziMainzicompute23 (gzdLLziMainzicompute23[130:67], gzdLLziMainzicompute23[66:3], gzdLLziMainzicompute23[2:0], callResR8);
  assign gzdLLziMainzicompute23R1 = {gzdLLziMainzicompute24[128:65], gzdLLziMainzicompute24[64:1], 3'h1};
  zdLLziMainzicompute23  zdLLziMainzicompute23R1 (gzdLLziMainzicompute23R1[130:67], gzdLLziMainzicompute23R1[66:3], gzdLLziMainzicompute23R1[2:0], callResR9);
  assign gzdLLziMainzicompute23R2 = {gzdLLziMainzicompute24[128:65], gzdLLziMainzicompute24[64:1], 3'h2};
  zdLLziMainzicompute23  zdLLziMainzicompute23R2 (gzdLLziMainzicompute23R2[130:67], gzdLLziMainzicompute23R2[66:3], gzdLLziMainzicompute23R2[2:0], callResR10);
  assign gzdLLziMainzicompute23R3 = {gzdLLziMainzicompute24[128:65], gzdLLziMainzicompute24[64:1], 3'h3};
  zdLLziMainzicompute23  zdLLziMainzicompute23R3 (gzdLLziMainzicompute23R3[130:67], gzdLLziMainzicompute23R3[66:3], gzdLLziMainzicompute23R3[2:0], callResR11);
  assign gzdLLziMainzicompute23R4 = {gzdLLziMainzicompute24[128:65], gzdLLziMainzicompute24[64:1], 3'h4};
  zdLLziMainzicompute23  zdLLziMainzicompute23R4 (gzdLLziMainzicompute23R4[130:67], gzdLLziMainzicompute23R4[66:3], gzdLLziMainzicompute23R4[2:0], callResR12);
  assign gzdLLziMainzicompute23R5 = {gzdLLziMainzicompute24[128:65], gzdLLziMainzicompute24[64:1], 3'h5};
  zdLLziMainzicompute23  zdLLziMainzicompute23R5 (gzdLLziMainzicompute23R5[130:67], gzdLLziMainzicompute23R5[66:3], gzdLLziMainzicompute23R5[2:0], callResR13);
  assign gzdLLziMainzicompute23R6 = {gzdLLziMainzicompute24[128:65], gzdLLziMainzicompute24[64:1], 3'h6};
  zdLLziMainzicompute23  zdLLziMainzicompute23R6 (gzdLLziMainzicompute23R6[130:67], gzdLLziMainzicompute23R6[66:3], gzdLLziMainzicompute23R6[2:0], callResR14);
  assign gzdLLziMainzicompute23R7 = {gzdLLziMainzicompute24[128:65], gzdLLziMainzicompute24[64:1], 3'h7};
  zdLLziMainzicompute23  zdLLziMainzicompute23R7 (gzdLLziMainzicompute23R7[130:67], gzdLLziMainzicompute23R7[66:3], gzdLLziMainzicompute23R7[2:0], callResR15);
  assign resizzeR9 = {callResR8, callResR9, callResR10, callResR11, callResR12, callResR13, callResR14, callResR15};
  assign resizzeR10 = gzdLLziMainzicompute24[131:129];
  assign binOpR10 = {128'(resizzeR10[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR11 = {binOpR10[255:128] * binOpR10[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR11 = binOpR11[255:128] % binOpR11[127:0];
  assign resizzeR12 = resizzeR11[2:0];
  assign binOpR12 = {128'h00000000000000000000000000000008, 128'(resizzeR12[2:0])};
  assign binOpR13 = {binOpR12[255:128] - binOpR12[127:0], 128'h00000000000000000000000000000001};
  assign binOpR14 = {binOpR13[255:128] - binOpR13[127:0], 128'h00000000000000000000000000000008};
  assign binOpR15 = {128'(resizzeR9[63:0]), binOpR14[255:128] * binOpR14[127:0]};
  assign resizzeR13 = binOpR15[255:128] >> binOpR15[127:0];
  assign res = (gzdLLziMainzicompute24[0] == 1'h1) ? resizzeR13[7:0] : resizzeR8[7:0];
endmodule

module zdLLziMainzicompute33 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [67:0] gzdLLziMainzicompute1;
  logic [7:0] callRes;
  logic [67:0] gzdLLziMainzicompute;
  logic [7:0] callResR1;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLziMainzicompute1 = {arg1, arg2, binOpR1[255:128] < binOpR1[127:0]};
  zdLLziMainzicompute1  zdLLziMainzicompute1 (gzdLLziMainzicompute1[67:4], gzdLLziMainzicompute1[3:1], callRes);
  assign gzdLLziMainzicompute = {arg0, arg2, binOp[255:128] < binOp[127:0]};
  zdLLziMainzicompute  zdLLziMainzicompute (gzdLLziMainzicompute[67:4], gzdLLziMainzicompute[3:1], callResR1);
  assign res = (gzdLLziMainzicompute[0] == 1'h1) ? callResR1 : callRes;
endmodule

module zdLLziMainzicompute37 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [67:0] gzdLLziMainzicompute15;
  logic [7:0] callRes;
  logic [67:0] gzdLLziMainzicompute14;
  logic [7:0] callResR1;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLziMainzicompute15 = {arg1, arg2, binOpR1[255:128] < binOpR1[127:0]};
  zdLLziMainzicompute15  zdLLziMainzicompute15 (gzdLLziMainzicompute15[67:4], gzdLLziMainzicompute15[3:1], callRes);
  assign gzdLLziMainzicompute14 = {arg0, arg2, binOp[255:128] < binOp[127:0]};
  zdLLziMainzicompute14  zdLLziMainzicompute14 (gzdLLziMainzicompute14[67:4], gzdLLziMainzicompute14[3:1], callResR1);
  assign res = (gzdLLziMainzicompute14[0] == 1'h1) ? callResR1 : callRes;
endmodule

module zdLLziMainzicompute39 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [255:0] binOp;
  logic [2:0] resizzeR1;
  logic [255:0] binOpR1;
  logic [131:0] gzdLLziMainzicompute38;
  logic [130:0] gzdLLziMainzicompute37;
  logic [7:0] callRes;
  logic [130:0] gzdLLziMainzicompute37R1;
  logic [7:0] callResR1;
  logic [130:0] gzdLLziMainzicompute37R2;
  logic [7:0] callResR2;
  logic [130:0] gzdLLziMainzicompute37R3;
  logic [7:0] callResR3;
  logic [130:0] gzdLLziMainzicompute37R4;
  logic [7:0] callResR4;
  logic [130:0] gzdLLziMainzicompute37R5;
  logic [7:0] callResR5;
  logic [130:0] gzdLLziMainzicompute37R6;
  logic [7:0] callResR6;
  logic [130:0] gzdLLziMainzicompute37R7;
  logic [7:0] callResR7;
  logic [63:0] resizzeR2;
  logic [2:0] resizzeR3;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR6;
  logic [2:0] resizzeR7;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [127:0] resizzeR8;
  logic [2:0] resizzeR9;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [127:0] resizzeR10;
  logic [131:0] gzdLLziMainzicompute34;
  logic [130:0] gzdLLziMainzicompute33;
  logic [7:0] callResR8;
  logic [130:0] gzdLLziMainzicompute33R1;
  logic [7:0] callResR9;
  logic [130:0] gzdLLziMainzicompute33R2;
  logic [7:0] callResR10;
  logic [130:0] gzdLLziMainzicompute33R3;
  logic [7:0] callResR11;
  logic [130:0] gzdLLziMainzicompute33R4;
  logic [7:0] callResR12;
  logic [130:0] gzdLLziMainzicompute33R5;
  logic [7:0] callResR13;
  logic [130:0] gzdLLziMainzicompute33R6;
  logic [7:0] callResR14;
  logic [130:0] gzdLLziMainzicompute33R7;
  logic [7:0] callResR15;
  logic [63:0] resizzeR11;
  logic [2:0] resizzeR12;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [127:0] resizzeR13;
  logic [2:0] resizzeR14;
  logic [255:0] binOpR14;
  logic [255:0] binOpR15;
  logic [127:0] resizzeR15;
  logic [2:0] resizzeR16;
  logic [255:0] binOpR16;
  logic [255:0] binOpR17;
  logic [255:0] binOpR18;
  logic [255:0] binOpR19;
  logic [127:0] resizzeR17;
  assign resizze = arg2;
  assign binOp = {128'(resizze[2:0]), 128'h00000000000000000000000000000003};
  assign resizzeR1 = arg2;
  assign binOpR1 = {128'(resizzeR1[2:0]), 128'h00000000000000000000000000000003};
  assign gzdLLziMainzicompute38 = {arg2, arg0, arg1, binOpR1[255:128] < binOpR1[127:0]};
  assign gzdLLziMainzicompute37 = {gzdLLziMainzicompute38[128:65], gzdLLziMainzicompute38[64:1], 3'h0};
  zdLLziMainzicompute37  zdLLziMainzicompute37 (gzdLLziMainzicompute37[130:67], gzdLLziMainzicompute37[66:3], gzdLLziMainzicompute37[2:0], callRes);
  assign gzdLLziMainzicompute37R1 = {gzdLLziMainzicompute38[128:65], gzdLLziMainzicompute38[64:1], 3'h1};
  zdLLziMainzicompute37  zdLLziMainzicompute37R1 (gzdLLziMainzicompute37R1[130:67], gzdLLziMainzicompute37R1[66:3], gzdLLziMainzicompute37R1[2:0], callResR1);
  assign gzdLLziMainzicompute37R2 = {gzdLLziMainzicompute38[128:65], gzdLLziMainzicompute38[64:1], 3'h2};
  zdLLziMainzicompute37  zdLLziMainzicompute37R2 (gzdLLziMainzicompute37R2[130:67], gzdLLziMainzicompute37R2[66:3], gzdLLziMainzicompute37R2[2:0], callResR2);
  assign gzdLLziMainzicompute37R3 = {gzdLLziMainzicompute38[128:65], gzdLLziMainzicompute38[64:1], 3'h3};
  zdLLziMainzicompute37  zdLLziMainzicompute37R3 (gzdLLziMainzicompute37R3[130:67], gzdLLziMainzicompute37R3[66:3], gzdLLziMainzicompute37R3[2:0], callResR3);
  assign gzdLLziMainzicompute37R4 = {gzdLLziMainzicompute38[128:65], gzdLLziMainzicompute38[64:1], 3'h4};
  zdLLziMainzicompute37  zdLLziMainzicompute37R4 (gzdLLziMainzicompute37R4[130:67], gzdLLziMainzicompute37R4[66:3], gzdLLziMainzicompute37R4[2:0], callResR4);
  assign gzdLLziMainzicompute37R5 = {gzdLLziMainzicompute38[128:65], gzdLLziMainzicompute38[64:1], 3'h5};
  zdLLziMainzicompute37  zdLLziMainzicompute37R5 (gzdLLziMainzicompute37R5[130:67], gzdLLziMainzicompute37R5[66:3], gzdLLziMainzicompute37R5[2:0], callResR5);
  assign gzdLLziMainzicompute37R6 = {gzdLLziMainzicompute38[128:65], gzdLLziMainzicompute38[64:1], 3'h6};
  zdLLziMainzicompute37  zdLLziMainzicompute37R6 (gzdLLziMainzicompute37R6[130:67], gzdLLziMainzicompute37R6[66:3], gzdLLziMainzicompute37R6[2:0], callResR6);
  assign gzdLLziMainzicompute37R7 = {gzdLLziMainzicompute38[128:65], gzdLLziMainzicompute38[64:1], 3'h7};
  zdLLziMainzicompute37  zdLLziMainzicompute37R7 (gzdLLziMainzicompute37R7[130:67], gzdLLziMainzicompute37R7[66:3], gzdLLziMainzicompute37R7[2:0], callResR7);
  assign resizzeR2 = {callRes, callResR1, callResR2, callResR3, callResR4, callResR5, callResR6, callResR7};
  assign resizzeR3 = gzdLLziMainzicompute38[131:129];
  assign binOpR2 = {128'(resizzeR3[2:0]), 128'h00000000000000000000000000000003};
  assign binOpR3 = {binOpR2[255:128] - binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR4 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR5 = resizzeR4[2:0];
  assign binOpR4 = {128'(resizzeR5[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR5 = {binOpR4[255:128] * binOpR4[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR6 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR7 = resizzeR6[2:0];
  assign binOpR6 = {128'(resizzeR7[2:0]), 128'h00000000000000000000000000000001};
  assign binOpR7 = {binOpR6[255:128] + binOpR6[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR8 = binOpR7[255:128] % binOpR7[127:0];
  assign resizzeR9 = resizzeR8[2:0];
  assign binOpR8 = {128'h00000000000000000000000000000008, 128'(resizzeR9[2:0])};
  assign binOpR9 = {binOpR8[255:128] - binOpR8[127:0], 128'h00000000000000000000000000000001};
  assign binOpR10 = {binOpR9[255:128] - binOpR9[127:0], 128'h00000000000000000000000000000008};
  assign binOpR11 = {128'(resizzeR2[63:0]), binOpR10[255:128] * binOpR10[127:0]};
  assign resizzeR10 = binOpR11[255:128] >> binOpR11[127:0];
  assign gzdLLziMainzicompute34 = {arg2, arg0, arg1, binOp[255:128] < binOp[127:0]};
  assign gzdLLziMainzicompute33 = {gzdLLziMainzicompute34[128:65], gzdLLziMainzicompute34[64:1], 3'h0};
  zdLLziMainzicompute33  zdLLziMainzicompute33 (gzdLLziMainzicompute33[130:67], gzdLLziMainzicompute33[66:3], gzdLLziMainzicompute33[2:0], callResR8);
  assign gzdLLziMainzicompute33R1 = {gzdLLziMainzicompute34[128:65], gzdLLziMainzicompute34[64:1], 3'h1};
  zdLLziMainzicompute33  zdLLziMainzicompute33R1 (gzdLLziMainzicompute33R1[130:67], gzdLLziMainzicompute33R1[66:3], gzdLLziMainzicompute33R1[2:0], callResR9);
  assign gzdLLziMainzicompute33R2 = {gzdLLziMainzicompute34[128:65], gzdLLziMainzicompute34[64:1], 3'h2};
  zdLLziMainzicompute33  zdLLziMainzicompute33R2 (gzdLLziMainzicompute33R2[130:67], gzdLLziMainzicompute33R2[66:3], gzdLLziMainzicompute33R2[2:0], callResR10);
  assign gzdLLziMainzicompute33R3 = {gzdLLziMainzicompute34[128:65], gzdLLziMainzicompute34[64:1], 3'h3};
  zdLLziMainzicompute33  zdLLziMainzicompute33R3 (gzdLLziMainzicompute33R3[130:67], gzdLLziMainzicompute33R3[66:3], gzdLLziMainzicompute33R3[2:0], callResR11);
  assign gzdLLziMainzicompute33R4 = {gzdLLziMainzicompute34[128:65], gzdLLziMainzicompute34[64:1], 3'h4};
  zdLLziMainzicompute33  zdLLziMainzicompute33R4 (gzdLLziMainzicompute33R4[130:67], gzdLLziMainzicompute33R4[66:3], gzdLLziMainzicompute33R4[2:0], callResR12);
  assign gzdLLziMainzicompute33R5 = {gzdLLziMainzicompute34[128:65], gzdLLziMainzicompute34[64:1], 3'h5};
  zdLLziMainzicompute33  zdLLziMainzicompute33R5 (gzdLLziMainzicompute33R5[130:67], gzdLLziMainzicompute33R5[66:3], gzdLLziMainzicompute33R5[2:0], callResR13);
  assign gzdLLziMainzicompute33R6 = {gzdLLziMainzicompute34[128:65], gzdLLziMainzicompute34[64:1], 3'h6};
  zdLLziMainzicompute33  zdLLziMainzicompute33R6 (gzdLLziMainzicompute33R6[130:67], gzdLLziMainzicompute33R6[66:3], gzdLLziMainzicompute33R6[2:0], callResR14);
  assign gzdLLziMainzicompute33R7 = {gzdLLziMainzicompute34[128:65], gzdLLziMainzicompute34[64:1], 3'h7};
  zdLLziMainzicompute33  zdLLziMainzicompute33R7 (gzdLLziMainzicompute33R7[130:67], gzdLLziMainzicompute33R7[66:3], gzdLLziMainzicompute33R7[2:0], callResR15);
  assign resizzeR11 = {callResR8, callResR9, callResR10, callResR11, callResR12, callResR13, callResR14, callResR15};
  assign resizzeR12 = gzdLLziMainzicompute34[131:129];
  assign binOpR12 = {128'(resizzeR12[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR13 = {binOpR12[255:128] * binOpR12[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR13 = binOpR13[255:128] % binOpR13[127:0];
  assign resizzeR14 = resizzeR13[2:0];
  assign binOpR14 = {128'(resizzeR14[2:0]), 128'h00000000000000000000000000000001};
  assign binOpR15 = {binOpR14[255:128] + binOpR14[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR15 = binOpR15[255:128] % binOpR15[127:0];
  assign resizzeR16 = resizzeR15[2:0];
  assign binOpR16 = {128'h00000000000000000000000000000008, 128'(resizzeR16[2:0])};
  assign binOpR17 = {binOpR16[255:128] - binOpR16[127:0], 128'h00000000000000000000000000000001};
  assign binOpR18 = {binOpR17[255:128] - binOpR17[127:0], 128'h00000000000000000000000000000008};
  assign binOpR19 = {128'(resizzeR11[63:0]), binOpR18[255:128] * binOpR18[127:0]};
  assign resizzeR17 = binOpR19[255:128] >> binOpR19[127:0];
  assign res = (gzdLLziMainzicompute34[0] == 1'h1) ? resizzeR17[7:0] : resizzeR10[7:0];
endmodule

module zdLLziMainzicompute41 (input logic [63:0] arg0,
  input logic [63:0] arg1,
  input logic [2:0] arg2,
  output logic [7:0] res);
  logic [2:0] resizze;
  logic [127:0] resizzeR1;
  logic [0:0] msbit;
  logic [0:0] gReWireziPreludezinot;
  logic [0:0] callRes;
  logic [2:0] resizzeR2;
  logic [127:0] resizzeR3;
  logic [0:0] msbitR1;
  logic [0:0] gReWireziPreludezinotR1;
  logic [0:0] callResR1;
  logic [131:0] gzdLLziMainzicompute40;
  logic [130:0] gzdLLziMainzicompute39;
  logic [7:0] callResR2;
  logic [130:0] gzdLLziMainzicompute39R1;
  logic [7:0] callResR3;
  logic [130:0] gzdLLziMainzicompute39R2;
  logic [7:0] callResR4;
  logic [130:0] gzdLLziMainzicompute39R3;
  logic [7:0] callResR5;
  logic [130:0] gzdLLziMainzicompute39R4;
  logic [7:0] callResR6;
  logic [130:0] gzdLLziMainzicompute39R5;
  logic [7:0] callResR7;
  logic [130:0] gzdLLziMainzicompute39R6;
  logic [7:0] callResR8;
  logic [130:0] gzdLLziMainzicompute39R7;
  logic [7:0] callResR9;
  logic [63:0] resizzeR4;
  logic [2:0] resizzeR5;
  logic [255:0] binOp;
  logic [255:0] binOpR1;
  logic [127:0] resizzeR6;
  logic [2:0] resizzeR7;
  logic [255:0] binOpR2;
  logic [255:0] binOpR3;
  logic [127:0] resizzeR8;
  logic [2:0] resizzeR9;
  logic [255:0] binOpR4;
  logic [255:0] binOpR5;
  logic [127:0] resizzeR10;
  logic [2:0] resizzeR11;
  logic [255:0] binOpR6;
  logic [255:0] binOpR7;
  logic [255:0] binOpR8;
  logic [255:0] binOpR9;
  logic [127:0] resizzeR12;
  logic [131:0] gzdLLziMainzicompute30;
  logic [130:0] gzdLLziMainzicompute29;
  logic [7:0] callResR10;
  logic [130:0] gzdLLziMainzicompute29R1;
  logic [7:0] callResR11;
  logic [130:0] gzdLLziMainzicompute29R2;
  logic [7:0] callResR12;
  logic [130:0] gzdLLziMainzicompute29R3;
  logic [7:0] callResR13;
  logic [130:0] gzdLLziMainzicompute29R4;
  logic [7:0] callResR14;
  logic [130:0] gzdLLziMainzicompute29R5;
  logic [7:0] callResR15;
  logic [130:0] gzdLLziMainzicompute29R6;
  logic [7:0] callResR16;
  logic [130:0] gzdLLziMainzicompute29R7;
  logic [7:0] callResR17;
  logic [63:0] resizzeR13;
  logic [2:0] resizzeR14;
  logic [255:0] binOpR10;
  logic [255:0] binOpR11;
  logic [127:0] resizzeR15;
  logic [2:0] resizzeR16;
  logic [255:0] binOpR12;
  logic [255:0] binOpR13;
  logic [127:0] resizzeR17;
  logic [2:0] resizzeR18;
  logic [255:0] binOpR14;
  logic [255:0] binOpR15;
  logic [255:0] binOpR16;
  logic [255:0] binOpR17;
  logic [127:0] resizzeR19;
  assign resizze = arg2;
  assign resizzeR1 = 128'(resizze[2:0]);
  assign msbit = resizzeR1[0];
  assign gReWireziPreludezinot = msbit[0];
  ReWireziPreludezinot  ReWireziPreludezinot (gReWireziPreludezinot[0], callRes);
  assign resizzeR2 = arg2;
  assign resizzeR3 = 128'(resizzeR2[2:0]);
  assign msbitR1 = resizzeR3[0];
  assign gReWireziPreludezinotR1 = msbitR1[0];
  ReWireziPreludezinot  ReWireziPreludezinotR1 (gReWireziPreludezinotR1[0], callResR1);
  assign gzdLLziMainzicompute40 = {arg0, arg1, arg2, callResR1};
  assign gzdLLziMainzicompute39 = {gzdLLziMainzicompute40[131:68], gzdLLziMainzicompute40[67:4], 3'h0};
  zdLLziMainzicompute39  zdLLziMainzicompute39 (gzdLLziMainzicompute39[130:67], gzdLLziMainzicompute39[66:3], gzdLLziMainzicompute39[2:0], callResR2);
  assign gzdLLziMainzicompute39R1 = {gzdLLziMainzicompute40[131:68], gzdLLziMainzicompute40[67:4], 3'h1};
  zdLLziMainzicompute39  zdLLziMainzicompute39R1 (gzdLLziMainzicompute39R1[130:67], gzdLLziMainzicompute39R1[66:3], gzdLLziMainzicompute39R1[2:0], callResR3);
  assign gzdLLziMainzicompute39R2 = {gzdLLziMainzicompute40[131:68], gzdLLziMainzicompute40[67:4], 3'h2};
  zdLLziMainzicompute39  zdLLziMainzicompute39R2 (gzdLLziMainzicompute39R2[130:67], gzdLLziMainzicompute39R2[66:3], gzdLLziMainzicompute39R2[2:0], callResR4);
  assign gzdLLziMainzicompute39R3 = {gzdLLziMainzicompute40[131:68], gzdLLziMainzicompute40[67:4], 3'h3};
  zdLLziMainzicompute39  zdLLziMainzicompute39R3 (gzdLLziMainzicompute39R3[130:67], gzdLLziMainzicompute39R3[66:3], gzdLLziMainzicompute39R3[2:0], callResR5);
  assign gzdLLziMainzicompute39R4 = {gzdLLziMainzicompute40[131:68], gzdLLziMainzicompute40[67:4], 3'h4};
  zdLLziMainzicompute39  zdLLziMainzicompute39R4 (gzdLLziMainzicompute39R4[130:67], gzdLLziMainzicompute39R4[66:3], gzdLLziMainzicompute39R4[2:0], callResR6);
  assign gzdLLziMainzicompute39R5 = {gzdLLziMainzicompute40[131:68], gzdLLziMainzicompute40[67:4], 3'h5};
  zdLLziMainzicompute39  zdLLziMainzicompute39R5 (gzdLLziMainzicompute39R5[130:67], gzdLLziMainzicompute39R5[66:3], gzdLLziMainzicompute39R5[2:0], callResR7);
  assign gzdLLziMainzicompute39R6 = {gzdLLziMainzicompute40[131:68], gzdLLziMainzicompute40[67:4], 3'h6};
  zdLLziMainzicompute39  zdLLziMainzicompute39R6 (gzdLLziMainzicompute39R6[130:67], gzdLLziMainzicompute39R6[66:3], gzdLLziMainzicompute39R6[2:0], callResR8);
  assign gzdLLziMainzicompute39R7 = {gzdLLziMainzicompute40[131:68], gzdLLziMainzicompute40[67:4], 3'h7};
  zdLLziMainzicompute39  zdLLziMainzicompute39R7 (gzdLLziMainzicompute39R7[130:67], gzdLLziMainzicompute39R7[66:3], gzdLLziMainzicompute39R7[2:0], callResR9);
  assign resizzeR4 = {callResR2, callResR3, callResR4, callResR5, callResR6, callResR7, callResR8, callResR9};
  assign resizzeR5 = gzdLLziMainzicompute40[3:1];
  assign binOp = {128'(resizzeR5[2:0]), 128'h00000000000000000000000000000001};
  assign binOpR1 = {binOp[255:128] - binOp[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR6 = binOpR1[255:128] % binOpR1[127:0];
  assign resizzeR7 = resizzeR6[2:0];
  assign binOpR2 = {128'h00000000000000000000000000000003, 128'(resizzeR7[2:0])};
  assign binOpR3 = {binOpR2[255:128] + binOpR2[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR8 = binOpR3[255:128] % binOpR3[127:0];
  assign resizzeR9 = resizzeR8[2:0];
  assign binOpR4 = {128'(resizzeR9[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR5 = {binOpR4[255:128] / binOpR4[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR10 = binOpR5[255:128] % binOpR5[127:0];
  assign resizzeR11 = resizzeR10[2:0];
  assign binOpR6 = {128'h00000000000000000000000000000008, 128'(resizzeR11[2:0])};
  assign binOpR7 = {binOpR6[255:128] - binOpR6[127:0], 128'h00000000000000000000000000000001};
  assign binOpR8 = {binOpR7[255:128] - binOpR7[127:0], 128'h00000000000000000000000000000008};
  assign binOpR9 = {128'(resizzeR4[63:0]), binOpR8[255:128] * binOpR8[127:0]};
  assign resizzeR12 = binOpR9[255:128] >> binOpR9[127:0];
  assign gzdLLziMainzicompute30 = {arg0, arg1, arg2, callRes};
  assign gzdLLziMainzicompute29 = {gzdLLziMainzicompute30[131:68], gzdLLziMainzicompute30[67:4], 3'h0};
  zdLLziMainzicompute29  zdLLziMainzicompute29 (gzdLLziMainzicompute29[130:67], gzdLLziMainzicompute29[66:3], gzdLLziMainzicompute29[2:0], callResR10);
  assign gzdLLziMainzicompute29R1 = {gzdLLziMainzicompute30[131:68], gzdLLziMainzicompute30[67:4], 3'h1};
  zdLLziMainzicompute29  zdLLziMainzicompute29R1 (gzdLLziMainzicompute29R1[130:67], gzdLLziMainzicompute29R1[66:3], gzdLLziMainzicompute29R1[2:0], callResR11);
  assign gzdLLziMainzicompute29R2 = {gzdLLziMainzicompute30[131:68], gzdLLziMainzicompute30[67:4], 3'h2};
  zdLLziMainzicompute29  zdLLziMainzicompute29R2 (gzdLLziMainzicompute29R2[130:67], gzdLLziMainzicompute29R2[66:3], gzdLLziMainzicompute29R2[2:0], callResR12);
  assign gzdLLziMainzicompute29R3 = {gzdLLziMainzicompute30[131:68], gzdLLziMainzicompute30[67:4], 3'h3};
  zdLLziMainzicompute29  zdLLziMainzicompute29R3 (gzdLLziMainzicompute29R3[130:67], gzdLLziMainzicompute29R3[66:3], gzdLLziMainzicompute29R3[2:0], callResR13);
  assign gzdLLziMainzicompute29R4 = {gzdLLziMainzicompute30[131:68], gzdLLziMainzicompute30[67:4], 3'h4};
  zdLLziMainzicompute29  zdLLziMainzicompute29R4 (gzdLLziMainzicompute29R4[130:67], gzdLLziMainzicompute29R4[66:3], gzdLLziMainzicompute29R4[2:0], callResR14);
  assign gzdLLziMainzicompute29R5 = {gzdLLziMainzicompute30[131:68], gzdLLziMainzicompute30[67:4], 3'h5};
  zdLLziMainzicompute29  zdLLziMainzicompute29R5 (gzdLLziMainzicompute29R5[130:67], gzdLLziMainzicompute29R5[66:3], gzdLLziMainzicompute29R5[2:0], callResR15);
  assign gzdLLziMainzicompute29R6 = {gzdLLziMainzicompute30[131:68], gzdLLziMainzicompute30[67:4], 3'h6};
  zdLLziMainzicompute29  zdLLziMainzicompute29R6 (gzdLLziMainzicompute29R6[130:67], gzdLLziMainzicompute29R6[66:3], gzdLLziMainzicompute29R6[2:0], callResR16);
  assign gzdLLziMainzicompute29R7 = {gzdLLziMainzicompute30[131:68], gzdLLziMainzicompute30[67:4], 3'h7};
  zdLLziMainzicompute29  zdLLziMainzicompute29R7 (gzdLLziMainzicompute29R7[130:67], gzdLLziMainzicompute29R7[66:3], gzdLLziMainzicompute29R7[2:0], callResR17);
  assign resizzeR13 = {callResR10, callResR11, callResR12, callResR13, callResR14, callResR15, callResR16, callResR17};
  assign resizzeR14 = gzdLLziMainzicompute30[3:1];
  assign binOpR10 = {128'h00000000000000000000000000000003, 128'(resizzeR14[2:0])};
  assign binOpR11 = {binOpR10[255:128] + binOpR10[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR15 = binOpR11[255:128] % binOpR11[127:0];
  assign resizzeR16 = resizzeR15[2:0];
  assign binOpR12 = {128'(resizzeR16[2:0]), 128'h00000000000000000000000000000002};
  assign binOpR13 = {binOpR12[255:128] / binOpR12[127:0], 128'h00000000000000000000000000000008};
  assign resizzeR17 = binOpR13[255:128] % binOpR13[127:0];
  assign resizzeR18 = resizzeR17[2:0];
  assign binOpR14 = {128'h00000000000000000000000000000008, 128'(resizzeR18[2:0])};
  assign binOpR15 = {binOpR14[255:128] - binOpR14[127:0], 128'h00000000000000000000000000000001};
  assign binOpR16 = {binOpR15[255:128] - binOpR15[127:0], 128'h00000000000000000000000000000008};
  assign binOpR17 = {128'(resizzeR13[63:0]), binOpR16[255:128] * binOpR16[127:0]};
  assign resizzeR19 = binOpR17[255:128] >> binOpR17[127:0];
  assign res = (gzdLLziMainzicompute30[0] == 1'h1) ? resizzeR19[7:0] : resizzeR12[7:0];
endmodule

module ReWireziPreludezinot (input logic [0:0] arg0,
  output logic [0:0] res);
  logic [0:0] lit;
  assign lit = arg0;
  assign res = (lit[0] == 1'h1) ? 1'h0 : 1'h1;
endmodule