module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [513:0] __in0,
  output logic [257:0] __out0);
  logic [1551:0] zll_pure_dispatch4_in;
  logic [1543:0] zll_pure_dispatch_in;
  logic [1543:0] zll_pure_dispatch14_in;
  logic [1543:0] zll_main_dev89_in;
  logic [1296:0] zll_main_dev89_out;
  logic [1551:0] zll_pure_dispatch16_in;
  logic [1543:0] zll_main_dev89_inR1;
  logic [1296:0] zll_main_dev89_outR1;
  logic [1551:0] zll_pure_dispatch8_in;
  logic [1543:0] zll_pure_dispatch9_in;
  logic [1543:0] zll_pure_dispatch11_in;
  logic [1543:0] zll_pure_dispatch7_in;
  logic [1543:0] main_dev_in;
  logic [1296:0] main_dev_out;
  logic [1551:0] zll_pure_dispatch6_in;
  logic [1549:0] zll_pure_dispatch10_in;
  logic [1549:0] zll_pure_dispatch3_in;
  logic [1549:0] zll_main_loop152_in;
  logic [1029:0] main_loop_in;
  logic [1296:0] main_loop_out;
  logic [1549:0] zll_main_loop125_in;
  logic [1543:0] zll_main_loop78_in;
  logic [1543:0] zll_main_loop88_in;
  logic [1285:0] zll_main_loop37_in;
  logic [1285:0] zll_main_loop145_in;
  logic [1285:0] zll_main_loop130_in;
  logic [1285:0] zll_main_loop85_in;
  logic [1285:0] zll_main_loop21_in;
  logic [1285:0] zll_main_loop143_in;
  logic [1285:0] zll_main_loop166_in;
  logic [1285:0] zll_main_loop47_in;
  logic [1285:0] zll_main_loop115_in;
  logic [1285:0] zll_main_loop135_in;
  logic [1285:0] zll_main_loop28_in;
  logic [1285:0] zll_main_loop161_in;
  logic [1285:0] zll_main_loop153_in;
  logic [1285:0] zll_main_loop118_in;
  logic [1285:0] zll_main_loop9_in;
  logic [1285:0] zll_main_loop105_in;
  logic [1285:0] zll_main_loop48_in;
  logic [1285:0] zll_main_loop43_in;
  logic [1541:0] zll_main_loop26_in;
  logic [1541:0] zll_main_loop138_in;
  logic [1541:0] zll_main_loop129_in;
  logic [1541:0] zll_main_loop24_in;
  logic [1541:0] zll_main_loop22_in;
  logic [1541:0] zll_main_loop127_in;
  logic [1541:0] zll_main_loop133_in;
  logic [1541:0] zll_main_loop100_in;
  logic [1541:0] zll_main_loop69_in;
  logic [1541:0] zll_main_loop68_in;
  logic [1541:0] zll_main_loop131_in;
  logic [1541:0] zll_main_loop59_in;
  logic [1541:0] zll_main_loop13_in;
  logic [1541:0] zll_main_loop120_in;
  logic [1541:0] zll_main_loop53_in;
  logic [1541:0] zll_main_loop25_in;
  logic [1541:0] zll_main_loop102_in;
  logic [1541:0] zll_main_loop155_in;
  logic [1541:0] zll_main_loop159_in;
  logic [1541:0] zll_main_loop110_in;
  logic [1541:0] zll_main_loop117_in;
  logic [1541:0] zll_main_loop90_in;
  logic [1541:0] zll_main_loop82_in;
  logic [1541:0] zll_main_loop99_in;
  logic [1541:0] zll_main_loop81_in;
  logic [1541:0] zll_main_loop139_in;
  logic [1541:0] zll_main_loop89_in;
  logic [1541:0] zll_main_loop98_in;
  logic [1541:0] zll_main_loop83_in;
  logic [63:0] plusw32_in;
  logic [31:0] extres;
  logic [63:0] plusw32_inR1;
  logic [31:0] extresR1;
  logic [63:0] plusw32_inR2;
  logic [31:0] extresR2;
  logic [63:0] plusw32_inR3;
  logic [31:0] extresR3;
  logic [63:0] plusw32_inR4;
  logic [31:0] extresR4;
  logic [63:0] plusw32_inR5;
  logic [31:0] extresR5;
  logic [63:0] plusw32_inR6;
  logic [31:0] extresR6;
  logic [63:0] plusw32_inR7;
  logic [31:0] extresR7;
  logic [1029:0] zll_main_loop16_in;
  logic [1029:0] zll_main_loop119_in;
  logic [1810:0] zll_main_loop70_in;
  logic [1810:0] zll_main_loop134_in;
  logic [1543:0] zll_main_loop114_in;
  logic [1543:0] zll_main_loop23_in;
  logic [1543:0] main_dev_inR1;
  logic [1296:0] main_dev_outR1;
  logic [0:0] __continue;
  logic [7:0] __resumption_tag;
  logic [223:0] __st0;
  logic [31:0] __st1;
  logic [511:0] __st2;
  logic [261:0] __st3;
  logic [7:0] __resumption_tag_next;
  logic [223:0] __st0_next;
  logic [31:0] __st1_next;
  logic [511:0] __st2_next;
  logic [261:0] __st3_next;
  assign zll_pure_dispatch4_in = {__in0, {__resumption_tag, __st0, __st1, __st2, __st3}};
  assign zll_pure_dispatch_in = {zll_pure_dispatch4_in[1551:1038], zll_pure_dispatch4_in[1029:774], zll_pure_dispatch4_in[773:262], zll_pure_dispatch4_in[261:6], zll_pure_dispatch4_in[5:0]};
  assign zll_pure_dispatch14_in = {zll_pure_dispatch_in[1029:774], zll_pure_dispatch_in[1543:1030], zll_pure_dispatch_in[773:262], zll_pure_dispatch_in[261:6], zll_pure_dispatch_in[5:0]};
  assign zll_main_dev89_in = {zll_pure_dispatch14_in[1287:774], zll_pure_dispatch14_in[1543:1288], zll_pure_dispatch14_in[773:262], zll_pure_dispatch14_in[261:6], zll_pure_dispatch14_in[5:0]};
  ZLL_Main_dev89  inst (zll_main_dev89_in[1543:1030], zll_main_dev89_in[1029:774], zll_main_dev89_in[773:262], zll_main_dev89_in[261:6], zll_main_dev89_in[5:0], zll_main_dev89_out);
  assign zll_pure_dispatch16_in = {__in0, {__resumption_tag, __st0, __st1, __st2, __st3}};
  assign zll_main_dev89_inR1 = {zll_pure_dispatch16_in[1551:1038], zll_pure_dispatch16_in[1029:774], zll_pure_dispatch16_in[773:262], zll_pure_dispatch16_in[261:6], zll_pure_dispatch16_in[5:0]};
  ZLL_Main_dev89  instR1 (zll_main_dev89_inR1[1543:1030], zll_main_dev89_inR1[1029:774], zll_main_dev89_inR1[773:262], zll_main_dev89_inR1[261:6], zll_main_dev89_inR1[5:0], zll_main_dev89_outR1);
  assign zll_pure_dispatch8_in = {__in0, {__resumption_tag, __st0, __st1, __st2, __st3}};
  assign zll_pure_dispatch9_in = {zll_pure_dispatch8_in[1551:1038], zll_pure_dispatch8_in[1029:774], zll_pure_dispatch8_in[773:262], zll_pure_dispatch8_in[261:6], zll_pure_dispatch8_in[5:0]};
  assign zll_pure_dispatch11_in = {zll_pure_dispatch9_in[1029:774], zll_pure_dispatch9_in[1543:1030], zll_pure_dispatch9_in[773:262], zll_pure_dispatch9_in[261:6], zll_pure_dispatch9_in[5:0]};
  assign zll_pure_dispatch7_in = {zll_pure_dispatch11_in[773:262], zll_pure_dispatch11_in[1543:1288], zll_pure_dispatch11_in[1287:774], zll_pure_dispatch11_in[261:6], zll_pure_dispatch11_in[5:0]};
  assign main_dev_in = {zll_pure_dispatch7_in[775:262], zll_pure_dispatch7_in[1031:776], zll_pure_dispatch7_in[1543:1032], zll_pure_dispatch7_in[261:6], zll_pure_dispatch7_in[5:0]};
  Main_dev  instR2 (main_dev_in[1543:1030], main_dev_in[1029:774], main_dev_in[773:262], main_dev_in[261:6], main_dev_in[5:0], main_dev_out);
  assign zll_pure_dispatch6_in = {__in0, {__resumption_tag, __st0, __st1, __st2, __st3}};
  assign zll_pure_dispatch10_in = {zll_pure_dispatch6_in[1551:1038], zll_pure_dispatch6_in[1035:1030], zll_pure_dispatch6_in[1029:774], zll_pure_dispatch6_in[773:262], zll_pure_dispatch6_in[261:6], zll_pure_dispatch6_in[5:0]};
  assign zll_pure_dispatch3_in = {zll_pure_dispatch10_in[1029:774], zll_pure_dispatch10_in[1549:1036], zll_pure_dispatch10_in[1035:1030], zll_pure_dispatch10_in[773:262], zll_pure_dispatch10_in[261:6], zll_pure_dispatch10_in[5:0]};
  assign zll_main_loop152_in = {zll_pure_dispatch3_in[779:774], zll_pure_dispatch3_in[1293:780], zll_pure_dispatch3_in[1549:1294], zll_pure_dispatch3_in[773:262], zll_pure_dispatch3_in[261:6], zll_pure_dispatch3_in[5:0]};
  assign main_loop_in = {zll_main_loop152_in[1029:774], zll_main_loop152_in[773:262], zll_main_loop152_in[261:6], zll_main_loop152_in[5:0]};
  Main_loop  instR3 (main_loop_in[1029:774], main_loop_in[773:262], main_loop_in[261:6], main_loop_in[5:0], main_loop_out);
  assign zll_main_loop125_in = {zll_main_loop152_in[5:0], zll_main_loop152_in[1029:774], zll_main_loop152_in[773:262], zll_main_loop152_in[261:6], zll_main_loop152_in[1543:1030], zll_main_loop152_in[1549:1544]};
  assign zll_main_loop78_in = {zll_main_loop125_in[1549:1544], zll_main_loop125_in[1543:1288], zll_main_loop125_in[1287:776], zll_main_loop125_in[775:520], zll_main_loop125_in[519:6]};
  assign zll_main_loop88_in = {zll_main_loop78_in[513:0], zll_main_loop78_in[1537:1282], zll_main_loop78_in[1281:770], zll_main_loop78_in[769:514], zll_main_loop78_in[1543:1538]};
  assign zll_main_loop37_in = {zll_main_loop88_in[261:6], zll_main_loop88_in[1029:774], zll_main_loop88_in[773:262], zll_main_loop88_in[261:6], zll_main_loop88_in[5:0]};
  assign zll_main_loop145_in = zll_main_loop37_in[1285:0];
  assign zll_main_loop130_in = {zll_main_loop145_in[1029:774], zll_main_loop145_in[1285:1030], zll_main_loop145_in[773:262], zll_main_loop145_in[261:6], zll_main_loop145_in[5:0]};
  assign zll_main_loop85_in = {zll_main_loop130_in[1285:1030], zll_main_loop130_in[773:262], zll_main_loop130_in[1029:774], zll_main_loop130_in[261:6], zll_main_loop130_in[5:0]};
  assign zll_main_loop21_in = {zll_main_loop85_in[517:262], zll_main_loop85_in[1285:1030], zll_main_loop85_in[1029:518], zll_main_loop85_in[261:6], zll_main_loop85_in[5:0]};
  assign zll_main_loop143_in = {zll_main_loop21_in[773:262], zll_main_loop21_in[5:0], zll_main_loop21_in[261:6], zll_main_loop21_in[1029:774], zll_main_loop21_in[1285:1030]};
  assign zll_main_loop166_in = {zll_main_loop143_in[1285:774], zll_main_loop143_in[255:224], zll_main_loop143_in[773:768], zll_main_loop143_in[767:512], zll_main_loop143_in[511:256], zll_main_loop143_in[223:192], zll_main_loop143_in[191:160], zll_main_loop143_in[159:128], zll_main_loop143_in[127:96], zll_main_loop143_in[95:64], zll_main_loop143_in[63:32], zll_main_loop143_in[31:0]};
  assign zll_main_loop47_in = {zll_main_loop166_in[1285:774], zll_main_loop166_in[773:742], zll_main_loop166_in[223:192], zll_main_loop166_in[741:736], zll_main_loop166_in[735:480], zll_main_loop166_in[479:224], zll_main_loop166_in[191:160], zll_main_loop166_in[159:128], zll_main_loop166_in[127:96], zll_main_loop166_in[95:64], zll_main_loop166_in[63:32], zll_main_loop166_in[31:0]};
  assign zll_main_loop115_in = {zll_main_loop47_in[1285:774], zll_main_loop47_in[191:160], zll_main_loop47_in[773:742], zll_main_loop47_in[741:710], zll_main_loop47_in[709:704], zll_main_loop47_in[703:448], zll_main_loop47_in[447:192], zll_main_loop47_in[159:128], zll_main_loop47_in[127:96], zll_main_loop47_in[95:64], zll_main_loop47_in[63:32], zll_main_loop47_in[31:0]};
  assign zll_main_loop135_in = {zll_main_loop115_in[1285:774], zll_main_loop115_in[159:128], zll_main_loop115_in[773:742], zll_main_loop115_in[741:710], zll_main_loop115_in[709:678], zll_main_loop115_in[677:672], zll_main_loop115_in[671:416], zll_main_loop115_in[415:160], zll_main_loop115_in[127:96], zll_main_loop115_in[95:64], zll_main_loop115_in[63:32], zll_main_loop115_in[31:0]};
  assign zll_main_loop28_in = {zll_main_loop135_in[1285:774], zll_main_loop135_in[773:742], zll_main_loop135_in[741:710], zll_main_loop135_in[709:678], zll_main_loop135_in[677:646], zll_main_loop135_in[127:96], zll_main_loop135_in[645:640], zll_main_loop135_in[639:384], zll_main_loop135_in[383:128], zll_main_loop135_in[95:64], zll_main_loop135_in[63:32], zll_main_loop135_in[31:0]};
  assign zll_main_loop161_in = {zll_main_loop28_in[1285:774], zll_main_loop28_in[773:742], zll_main_loop28_in[741:710], zll_main_loop28_in[709:678], zll_main_loop28_in[677:646], zll_main_loop28_in[645:614], zll_main_loop28_in[95:64], zll_main_loop28_in[613:608], zll_main_loop28_in[607:352], zll_main_loop28_in[351:96], zll_main_loop28_in[63:32], zll_main_loop28_in[31:0]};
  assign zll_main_loop153_in = {zll_main_loop161_in[1285:774], zll_main_loop161_in[773:742], zll_main_loop161_in[63:32], zll_main_loop161_in[741:710], zll_main_loop161_in[709:678], zll_main_loop161_in[677:646], zll_main_loop161_in[645:614], zll_main_loop161_in[613:582], zll_main_loop161_in[581:576], zll_main_loop161_in[575:320], zll_main_loop161_in[319:64], zll_main_loop161_in[31:0]};
  assign zll_main_loop118_in = {zll_main_loop153_in[677:646], zll_main_loop153_in[645:614], zll_main_loop153_in[709:678], zll_main_loop153_in[773:742], zll_main_loop153_in[613:582], zll_main_loop153_in[581:550], zll_main_loop153_in[741:710], zll_main_loop153_in[31:0], zll_main_loop153_in[287:32], zll_main_loop153_in[1285:774], zll_main_loop153_in[543:288], zll_main_loop153_in[549:544]};
  assign zll_main_loop9_in = {zll_main_loop118_in[1285:1254], zll_main_loop118_in[1221:1190], zll_main_loop118_in[1253:1222], zll_main_loop118_in[1189:1158], zll_main_loop118_in[1157:1126], zll_main_loop118_in[1125:1094], zll_main_loop118_in[1093:1062], zll_main_loop118_in[1061:1030], zll_main_loop118_in[1029:774], zll_main_loop118_in[773:262], zll_main_loop118_in[261:6], zll_main_loop118_in[5:0]};
  assign zll_main_loop105_in = {zll_main_loop9_in[1285:1254], zll_main_loop9_in[1253:1222], zll_main_loop9_in[1157:1126], zll_main_loop9_in[1221:1190], zll_main_loop9_in[1189:1158], zll_main_loop9_in[1125:1094], zll_main_loop9_in[1093:1062], zll_main_loop9_in[1061:1030], zll_main_loop9_in[1029:774], zll_main_loop9_in[773:262], zll_main_loop9_in[261:6], zll_main_loop9_in[5:0]};
  assign zll_main_loop48_in = {zll_main_loop105_in[1285:1254], zll_main_loop105_in[1253:1222], zll_main_loop105_in[1221:1190], zll_main_loop105_in[1125:1094], zll_main_loop105_in[1189:1158], zll_main_loop105_in[1157:1126], zll_main_loop105_in[1093:1062], zll_main_loop105_in[1061:1030], zll_main_loop105_in[1029:774], zll_main_loop105_in[773:262], zll_main_loop105_in[261:6], zll_main_loop105_in[5:0]};
  assign zll_main_loop43_in = {zll_main_loop48_in[1093:1062], zll_main_loop48_in[1285:1254], zll_main_loop48_in[1253:1222], zll_main_loop48_in[1221:1190], zll_main_loop48_in[1189:1158], zll_main_loop48_in[1157:1126], zll_main_loop48_in[1125:1094], zll_main_loop48_in[1061:1030], zll_main_loop48_in[1029:774], zll_main_loop48_in[773:262], zll_main_loop48_in[261:6], zll_main_loop48_in[5:0]};
  assign zll_main_loop26_in = {zll_main_loop43_in[1061:1030], zll_main_loop43_in[1125:1094], zll_main_loop43_in[1253:1222], zll_main_loop43_in[1093:1062], zll_main_loop43_in[1189:1158], zll_main_loop43_in[1221:1190], zll_main_loop43_in[1285:1254], zll_main_loop43_in[1157:1126], zll_main_loop43_in[1029:774], zll_main_loop43_in[1029:774], zll_main_loop43_in[773:262], zll_main_loop43_in[261:6], zll_main_loop43_in[5:0]};
  assign zll_main_loop138_in = {zll_main_loop26_in[1541:1510], zll_main_loop26_in[1509:1478], zll_main_loop26_in[1477:1446], zll_main_loop26_in[1445:1414], zll_main_loop26_in[1413:1382], zll_main_loop26_in[1381:1350], zll_main_loop26_in[1349:1318], zll_main_loop26_in[1317:1286], zll_main_loop26_in[1285:0]};
  assign zll_main_loop129_in = {zll_main_loop138_in[1541:1510], zll_main_loop138_in[1509:1478], zll_main_loop138_in[1477:1446], zll_main_loop138_in[1445:1414], zll_main_loop138_in[1413:1382], zll_main_loop138_in[1381:1350], zll_main_loop138_in[1349:1318], zll_main_loop138_in[1285:1030], zll_main_loop138_in[1317:1286], zll_main_loop138_in[1029:774], zll_main_loop138_in[773:262], zll_main_loop138_in[261:6], zll_main_loop138_in[5:0]};
  assign zll_main_loop24_in = {zll_main_loop129_in[1541:1510], zll_main_loop129_in[1509:1478], zll_main_loop129_in[1477:1446], zll_main_loop129_in[1445:1414], zll_main_loop129_in[1413:1382], zll_main_loop129_in[1381:1350], zll_main_loop129_in[1349:1318], zll_main_loop129_in[1029:774], zll_main_loop129_in[1317:1062], zll_main_loop129_in[1061:1030], zll_main_loop129_in[773:262], zll_main_loop129_in[261:6], zll_main_loop129_in[5:0]};
  assign zll_main_loop22_in = {zll_main_loop24_in[1541:1510], zll_main_loop24_in[1509:1478], zll_main_loop24_in[1477:1446], zll_main_loop24_in[1445:1414], zll_main_loop24_in[1413:1382], zll_main_loop24_in[1381:1350], zll_main_loop24_in[1349:1318], zll_main_loop24_in[1317:1062], zll_main_loop24_in[773:262], zll_main_loop24_in[1061:806], zll_main_loop24_in[805:774], zll_main_loop24_in[261:6], zll_main_loop24_in[5:0]};
  assign zll_main_loop127_in = {zll_main_loop22_in[1477:1446], zll_main_loop22_in[1349:1318], zll_main_loop22_in[293:262], zll_main_loop22_in[1413:1382], zll_main_loop22_in[1445:1414], zll_main_loop22_in[1541:1510], zll_main_loop22_in[1381:1350], zll_main_loop22_in[1509:1478], zll_main_loop22_in[549:294], zll_main_loop22_in[1317:1062], zll_main_loop22_in[1061:550], zll_main_loop22_in[261:6], zll_main_loop22_in[5:0]};
  assign zll_main_loop133_in = {zll_main_loop127_in[261:6], zll_main_loop127_in[1029:774], zll_main_loop127_in[773:262], zll_main_loop127_in[5:0], zll_main_loop127_in[1541:1510], zll_main_loop127_in[1445:1414], zll_main_loop127_in[1381:1350], zll_main_loop127_in[1477:1446], zll_main_loop127_in[1349:1318], zll_main_loop127_in[1509:1478], zll_main_loop127_in[1413:1382], zll_main_loop127_in[1317:1286], zll_main_loop127_in[1285:1030]};
  assign zll_main_loop100_in = {zll_main_loop133_in[1541:1286], zll_main_loop133_in[511:480], zll_main_loop133_in[1285:1030], zll_main_loop133_in[1029:518], zll_main_loop133_in[517:512], zll_main_loop133_in[479:448], zll_main_loop133_in[447:416], zll_main_loop133_in[415:384], zll_main_loop133_in[383:352], zll_main_loop133_in[351:320], zll_main_loop133_in[319:288], zll_main_loop133_in[287:256], zll_main_loop133_in[255:224], zll_main_loop133_in[223:192], zll_main_loop133_in[191:160], zll_main_loop133_in[159:128], zll_main_loop133_in[127:96], zll_main_loop133_in[95:64], zll_main_loop133_in[63:32], zll_main_loop133_in[31:0]};
  assign zll_main_loop69_in = {zll_main_loop100_in[1541:1286], zll_main_loop100_in[1285:1254], zll_main_loop100_in[1253:998], zll_main_loop100_in[479:448], zll_main_loop100_in[997:486], zll_main_loop100_in[485:480], zll_main_loop100_in[447:416], zll_main_loop100_in[415:384], zll_main_loop100_in[383:352], zll_main_loop100_in[351:320], zll_main_loop100_in[319:288], zll_main_loop100_in[287:256], zll_main_loop100_in[255:224], zll_main_loop100_in[223:192], zll_main_loop100_in[191:160], zll_main_loop100_in[159:128], zll_main_loop100_in[127:96], zll_main_loop100_in[95:64], zll_main_loop100_in[63:32], zll_main_loop100_in[31:0]};
  assign zll_main_loop68_in = {zll_main_loop69_in[1541:1286], zll_main_loop69_in[447:416], zll_main_loop69_in[1285:1254], zll_main_loop69_in[1253:998], zll_main_loop69_in[997:966], zll_main_loop69_in[965:454], zll_main_loop69_in[453:448], zll_main_loop69_in[415:384], zll_main_loop69_in[383:352], zll_main_loop69_in[351:320], zll_main_loop69_in[319:288], zll_main_loop69_in[287:256], zll_main_loop69_in[255:224], zll_main_loop69_in[223:192], zll_main_loop69_in[191:160], zll_main_loop69_in[159:128], zll_main_loop69_in[127:96], zll_main_loop69_in[95:64], zll_main_loop69_in[63:32], zll_main_loop69_in[31:0]};
  assign zll_main_loop131_in = {zll_main_loop68_in[1541:1286], zll_main_loop68_in[1285:1254], zll_main_loop68_in[1253:1222], zll_main_loop68_in[1221:966], zll_main_loop68_in[965:934], zll_main_loop68_in[933:422], zll_main_loop68_in[421:416], zll_main_loop68_in[383:352], zll_main_loop68_in[415:384], zll_main_loop68_in[351:320], zll_main_loop68_in[319:288], zll_main_loop68_in[287:256], zll_main_loop68_in[255:224], zll_main_loop68_in[223:192], zll_main_loop68_in[191:160], zll_main_loop68_in[159:128], zll_main_loop68_in[127:96], zll_main_loop68_in[95:64], zll_main_loop68_in[63:32], zll_main_loop68_in[31:0]};
  assign zll_main_loop59_in = {zll_main_loop131_in[1541:1286], zll_main_loop131_in[1285:1254], zll_main_loop131_in[1253:1222], zll_main_loop131_in[1221:966], zll_main_loop131_in[965:934], zll_main_loop131_in[933:422], zll_main_loop131_in[351:320], zll_main_loop131_in[421:416], zll_main_loop131_in[415:384], zll_main_loop131_in[383:352], zll_main_loop131_in[319:288], zll_main_loop131_in[287:256], zll_main_loop131_in[255:224], zll_main_loop131_in[223:192], zll_main_loop131_in[191:160], zll_main_loop131_in[159:128], zll_main_loop131_in[127:96], zll_main_loop131_in[95:64], zll_main_loop131_in[63:32], zll_main_loop131_in[31:0]};
  assign zll_main_loop13_in = {zll_main_loop59_in[1541:1286], zll_main_loop59_in[1285:1254], zll_main_loop59_in[1253:1222], zll_main_loop59_in[1221:966], zll_main_loop59_in[965:934], zll_main_loop59_in[933:422], zll_main_loop59_in[421:390], zll_main_loop59_in[319:288], zll_main_loop59_in[389:384], zll_main_loop59_in[383:352], zll_main_loop59_in[351:320], zll_main_loop59_in[287:256], zll_main_loop59_in[255:224], zll_main_loop59_in[223:192], zll_main_loop59_in[191:160], zll_main_loop59_in[159:128], zll_main_loop59_in[127:96], zll_main_loop59_in[95:64], zll_main_loop59_in[63:32], zll_main_loop59_in[31:0]};
  assign zll_main_loop120_in = {zll_main_loop13_in[1541:1286], zll_main_loop13_in[1285:1254], zll_main_loop13_in[287:256], zll_main_loop13_in[1253:1222], zll_main_loop13_in[1221:966], zll_main_loop13_in[965:934], zll_main_loop13_in[933:422], zll_main_loop13_in[421:390], zll_main_loop13_in[389:358], zll_main_loop13_in[357:352], zll_main_loop13_in[351:320], zll_main_loop13_in[319:288], zll_main_loop13_in[255:224], zll_main_loop13_in[223:192], zll_main_loop13_in[191:160], zll_main_loop13_in[159:128], zll_main_loop13_in[127:96], zll_main_loop13_in[95:64], zll_main_loop13_in[63:32], zll_main_loop13_in[31:0]};
  assign zll_main_loop53_in = {zll_main_loop120_in[1541:1286], zll_main_loop120_in[255:224], zll_main_loop120_in[1285:1254], zll_main_loop120_in[1253:1222], zll_main_loop120_in[1221:1190], zll_main_loop120_in[1189:934], zll_main_loop120_in[933:902], zll_main_loop120_in[901:390], zll_main_loop120_in[389:358], zll_main_loop120_in[357:326], zll_main_loop120_in[325:320], zll_main_loop120_in[319:288], zll_main_loop120_in[287:256], zll_main_loop120_in[223:192], zll_main_loop120_in[191:160], zll_main_loop120_in[159:128], zll_main_loop120_in[127:96], zll_main_loop120_in[95:64], zll_main_loop120_in[63:32], zll_main_loop120_in[31:0]};
  assign zll_main_loop25_in = {zll_main_loop53_in[1541:1286], zll_main_loop53_in[1285:1254], zll_main_loop53_in[1253:1222], zll_main_loop53_in[1221:1190], zll_main_loop53_in[1189:1158], zll_main_loop53_in[1157:902], zll_main_loop53_in[901:870], zll_main_loop53_in[223:192], zll_main_loop53_in[869:358], zll_main_loop53_in[357:326], zll_main_loop53_in[325:294], zll_main_loop53_in[293:288], zll_main_loop53_in[287:256], zll_main_loop53_in[255:224], zll_main_loop53_in[191:160], zll_main_loop53_in[159:128], zll_main_loop53_in[127:96], zll_main_loop53_in[95:64], zll_main_loop53_in[63:32], zll_main_loop53_in[31:0]};
  assign zll_main_loop102_in = {zll_main_loop25_in[1541:1286], zll_main_loop25_in[1285:1254], zll_main_loop25_in[1253:1222], zll_main_loop25_in[1221:1190], zll_main_loop25_in[1189:1158], zll_main_loop25_in[1157:902], zll_main_loop25_in[901:870], zll_main_loop25_in[869:838], zll_main_loop25_in[837:326], zll_main_loop25_in[325:294], zll_main_loop25_in[293:262], zll_main_loop25_in[191:160], zll_main_loop25_in[261:256], zll_main_loop25_in[255:224], zll_main_loop25_in[223:192], zll_main_loop25_in[159:128], zll_main_loop25_in[127:96], zll_main_loop25_in[95:64], zll_main_loop25_in[63:32], zll_main_loop25_in[31:0]};
  assign zll_main_loop155_in = {zll_main_loop102_in[1541:1286], zll_main_loop102_in[1285:1254], zll_main_loop102_in[1253:1222], zll_main_loop102_in[1221:1190], zll_main_loop102_in[1189:1158], zll_main_loop102_in[1157:902], zll_main_loop102_in[901:870], zll_main_loop102_in[869:838], zll_main_loop102_in[837:326], zll_main_loop102_in[325:294], zll_main_loop102_in[293:262], zll_main_loop102_in[261:230], zll_main_loop102_in[229:224], zll_main_loop102_in[159:128], zll_main_loop102_in[223:192], zll_main_loop102_in[191:160], zll_main_loop102_in[127:96], zll_main_loop102_in[95:64], zll_main_loop102_in[63:32], zll_main_loop102_in[31:0]};
  assign zll_main_loop159_in = {zll_main_loop155_in[1541:1286], zll_main_loop155_in[1285:1254], zll_main_loop155_in[1253:1222], zll_main_loop155_in[1221:1190], zll_main_loop155_in[1189:1158], zll_main_loop155_in[1157:902], zll_main_loop155_in[901:870], zll_main_loop155_in[869:838], zll_main_loop155_in[127:96], zll_main_loop155_in[837:326], zll_main_loop155_in[325:294], zll_main_loop155_in[293:262], zll_main_loop155_in[261:230], zll_main_loop155_in[229:224], zll_main_loop155_in[223:192], zll_main_loop155_in[191:160], zll_main_loop155_in[159:128], zll_main_loop155_in[95:64], zll_main_loop155_in[63:32], zll_main_loop155_in[31:0]};
  assign zll_main_loop110_in = {zll_main_loop159_in[1541:1286], zll_main_loop159_in[1285:1254], zll_main_loop159_in[1253:1222], zll_main_loop159_in[1221:1190], zll_main_loop159_in[1189:1158], zll_main_loop159_in[1157:902], zll_main_loop159_in[901:870], zll_main_loop159_in[869:838], zll_main_loop159_in[837:806], zll_main_loop159_in[805:294], zll_main_loop159_in[293:262], zll_main_loop159_in[261:230], zll_main_loop159_in[229:198], zll_main_loop159_in[197:192], zll_main_loop159_in[95:64], zll_main_loop159_in[191:160], zll_main_loop159_in[159:128], zll_main_loop159_in[127:96], zll_main_loop159_in[63:32], zll_main_loop159_in[31:0]};
  assign zll_main_loop117_in = {zll_main_loop110_in[1541:1286], zll_main_loop110_in[1285:1254], zll_main_loop110_in[1253:1222], zll_main_loop110_in[1221:1190], zll_main_loop110_in[1189:1158], zll_main_loop110_in[63:32], zll_main_loop110_in[1157:902], zll_main_loop110_in[901:870], zll_main_loop110_in[869:838], zll_main_loop110_in[837:806], zll_main_loop110_in[805:294], zll_main_loop110_in[293:262], zll_main_loop110_in[261:230], zll_main_loop110_in[229:198], zll_main_loop110_in[197:192], zll_main_loop110_in[191:160], zll_main_loop110_in[159:128], zll_main_loop110_in[127:96], zll_main_loop110_in[95:64], zll_main_loop110_in[31:0]};
  assign zll_main_loop90_in = {zll_main_loop117_in[1189:1158], zll_main_loop117_in[869:838], zll_main_loop117_in[1253:1222], zll_main_loop117_in[63:32], zll_main_loop117_in[95:64], zll_main_loop117_in[261:230], zll_main_loop117_in[229:198], zll_main_loop117_in[1221:1190], zll_main_loop117_in[1285:1254], zll_main_loop117_in[837:806], zll_main_loop117_in[197:166], zll_main_loop117_in[127:96], zll_main_loop117_in[805:774], zll_main_loop117_in[159:128], zll_main_loop117_in[1157:1126], zll_main_loop117_in[31:0], zll_main_loop117_in[1125:870], zll_main_loop117_in[773:262], zll_main_loop117_in[1541:1286], zll_main_loop117_in[165:160]};
  assign zll_main_loop82_in = {zll_main_loop90_in[1541:1510], zll_main_loop90_in[1509:1478], zll_main_loop90_in[1477:1446], zll_main_loop90_in[1445:1414], zll_main_loop90_in[1285:1254], zll_main_loop90_in[1413:1382], zll_main_loop90_in[1381:1350], zll_main_loop90_in[1349:1318], zll_main_loop90_in[1317:1286], zll_main_loop90_in[1253:1222], zll_main_loop90_in[1221:1190], zll_main_loop90_in[1189:1158], zll_main_loop90_in[1157:1126], zll_main_loop90_in[1125:1094], zll_main_loop90_in[1093:1062], zll_main_loop90_in[1061:1030], zll_main_loop90_in[1029:774], zll_main_loop90_in[773:262], zll_main_loop90_in[261:6], zll_main_loop90_in[5:0]};
  assign zll_main_loop99_in = {zll_main_loop82_in[1541:1510], zll_main_loop82_in[1509:1478], zll_main_loop82_in[1477:1446], zll_main_loop82_in[1253:1222], zll_main_loop82_in[1445:1414], zll_main_loop82_in[1413:1382], zll_main_loop82_in[1381:1350], zll_main_loop82_in[1349:1318], zll_main_loop82_in[1317:1286], zll_main_loop82_in[1285:1254], zll_main_loop82_in[1221:1190], zll_main_loop82_in[1189:1158], zll_main_loop82_in[1157:1126], zll_main_loop82_in[1125:1094], zll_main_loop82_in[1093:1062], zll_main_loop82_in[1061:1030], zll_main_loop82_in[1029:774], zll_main_loop82_in[773:262], zll_main_loop82_in[261:6], zll_main_loop82_in[5:0]};
  assign zll_main_loop81_in = {zll_main_loop99_in[1541:1510], zll_main_loop99_in[1509:1478], zll_main_loop99_in[1477:1446], zll_main_loop99_in[1445:1414], zll_main_loop99_in[1413:1382], zll_main_loop99_in[1381:1350], zll_main_loop99_in[1349:1318], zll_main_loop99_in[1221:1190], zll_main_loop99_in[1317:1286], zll_main_loop99_in[1285:1254], zll_main_loop99_in[1253:1222], zll_main_loop99_in[1189:1158], zll_main_loop99_in[1157:1126], zll_main_loop99_in[1125:1094], zll_main_loop99_in[1093:1062], zll_main_loop99_in[1061:1030], zll_main_loop99_in[1029:774], zll_main_loop99_in[773:262], zll_main_loop99_in[261:6], zll_main_loop99_in[5:0]};
  assign zll_main_loop139_in = {zll_main_loop81_in[1541:1510], zll_main_loop81_in[1509:1478], zll_main_loop81_in[1477:1446], zll_main_loop81_in[1445:1414], zll_main_loop81_in[1413:1382], zll_main_loop81_in[1189:1158], zll_main_loop81_in[1381:1350], zll_main_loop81_in[1349:1318], zll_main_loop81_in[1317:1286], zll_main_loop81_in[1285:1254], zll_main_loop81_in[1253:1222], zll_main_loop81_in[1221:1190], zll_main_loop81_in[1157:1126], zll_main_loop81_in[1125:1094], zll_main_loop81_in[1093:1062], zll_main_loop81_in[1061:1030], zll_main_loop81_in[1029:774], zll_main_loop81_in[773:262], zll_main_loop81_in[261:6], zll_main_loop81_in[5:0]};
  assign zll_main_loop89_in = {zll_main_loop139_in[1541:1510], zll_main_loop139_in[1509:1478], zll_main_loop139_in[1477:1446], zll_main_loop139_in[1445:1414], zll_main_loop139_in[1413:1382], zll_main_loop139_in[1381:1350], zll_main_loop139_in[1349:1318], zll_main_loop139_in[1317:1286], zll_main_loop139_in[1285:1254], zll_main_loop139_in[1157:1126], zll_main_loop139_in[1253:1222], zll_main_loop139_in[1221:1190], zll_main_loop139_in[1189:1158], zll_main_loop139_in[1125:1094], zll_main_loop139_in[1093:1062], zll_main_loop139_in[1061:1030], zll_main_loop139_in[1029:774], zll_main_loop139_in[773:262], zll_main_loop139_in[261:6], zll_main_loop139_in[5:0]};
  assign zll_main_loop98_in = {zll_main_loop89_in[1541:1510], zll_main_loop89_in[1509:1478], zll_main_loop89_in[1477:1446], zll_main_loop89_in[1125:1094], zll_main_loop89_in[1445:1414], zll_main_loop89_in[1413:1382], zll_main_loop89_in[1381:1350], zll_main_loop89_in[1349:1318], zll_main_loop89_in[1317:1286], zll_main_loop89_in[1285:1254], zll_main_loop89_in[1253:1222], zll_main_loop89_in[1221:1190], zll_main_loop89_in[1189:1158], zll_main_loop89_in[1157:1126], zll_main_loop89_in[1093:1062], zll_main_loop89_in[1061:1030], zll_main_loop89_in[1029:774], zll_main_loop89_in[773:262], zll_main_loop89_in[261:6], zll_main_loop89_in[5:0]};
  assign zll_main_loop83_in = {zll_main_loop98_in[1541:1510], zll_main_loop98_in[1509:1478], zll_main_loop98_in[1477:1446], zll_main_loop98_in[1445:1414], zll_main_loop98_in[1413:1382], zll_main_loop98_in[1381:1350], zll_main_loop98_in[1349:1318], zll_main_loop98_in[1317:1286], zll_main_loop98_in[1285:1254], zll_main_loop98_in[1253:1222], zll_main_loop98_in[1221:1190], zll_main_loop98_in[1189:1158], zll_main_loop98_in[1093:1062], zll_main_loop98_in[1157:1126], zll_main_loop98_in[1125:1094], zll_main_loop98_in[1061:1030], zll_main_loop98_in[1029:774], zll_main_loop98_in[773:262], zll_main_loop98_in[261:6], zll_main_loop98_in[5:0]};
  assign plusw32_in = {zll_main_loop83_in[1317:1286], zll_main_loop83_in[1541:1510]};
  plusW32  instR4 (plusw32_in[63:32], plusw32_in[31:0], extres[31:0]);
  assign plusw32_inR1 = {zll_main_loop83_in[1413:1382], zll_main_loop83_in[1093:1062]};
  plusW32  instR5 (plusw32_inR1[63:32], plusw32_inR1[31:0], extresR1[31:0]);
  assign plusw32_inR2 = {zll_main_loop83_in[1253:1222], zll_main_loop83_in[1285:1254]};
  plusW32  instR6 (plusw32_inR2[63:32], plusw32_inR2[31:0], extresR2[31:0]);
  assign plusw32_inR3 = {zll_main_loop83_in[1349:1318], zll_main_loop83_in[1125:1094]};
  plusW32  instR7 (plusw32_inR3[63:32], plusw32_inR3[31:0], extresR3[31:0]);
  assign plusw32_inR4 = {zll_main_loop83_in[1221:1190], zll_main_loop83_in[1509:1478]};
  plusW32  instR8 (plusw32_inR4[63:32], plusw32_inR4[31:0], extresR4[31:0]);
  assign plusw32_inR5 = {zll_main_loop83_in[1445:1414], zll_main_loop83_in[1381:1350]};
  plusW32  instR9 (plusw32_inR5[63:32], plusw32_inR5[31:0], extresR5[31:0]);
  assign plusw32_inR6 = {zll_main_loop83_in[1157:1126], zll_main_loop83_in[1189:1158]};
  plusW32  instR10 (plusw32_inR6[63:32], plusw32_inR6[31:0], extresR6[31:0]);
  assign plusw32_inR7 = {zll_main_loop83_in[1061:1030], zll_main_loop83_in[1477:1446]};
  plusW32  instR11 (plusw32_inR7[63:32], plusw32_inR7[31:0], extresR7[31:0]);
  assign zll_main_loop16_in = {zll_main_loop83_in[1029:774], zll_main_loop83_in[773:262], extres, extresR1, extresR2, extresR3, extresR4, extresR5, extresR6, extresR7, zll_main_loop83_in[5:0]};
  assign zll_main_loop119_in = zll_main_loop16_in[1029:0];
  assign zll_main_loop70_in = {zll_main_loop88_in[1543:1030], {{10'h1, {9'h101{1'h0}}}, zll_main_loop119_in[1029:774], zll_main_loop119_in[773:262], zll_main_loop119_in[261:6], zll_main_loop119_in[5:0]}};
  assign zll_main_loop134_in = {zll_main_loop70_in[1810:1297], zll_main_loop70_in[1296:0]};
  assign zll_main_loop114_in = {zll_main_loop134_in[1810:1297], zll_main_loop134_in[1029:774], zll_main_loop134_in[773:262], zll_main_loop134_in[261:6], zll_main_loop134_in[5:0]};
  assign zll_main_loop23_in = {zll_main_loop114_in[1543:1030], zll_main_loop114_in[773:262], zll_main_loop114_in[1029:774], zll_main_loop114_in[261:6], zll_main_loop114_in[5:0]};
  assign main_dev_inR1 = {zll_main_loop23_in[1543:1030], zll_main_loop23_in[517:262], zll_main_loop23_in[1029:518], zll_main_loop23_in[261:6], zll_main_loop23_in[5:0]};
  Main_dev  instR12 (main_dev_inR1[1543:1030], main_dev_inR1[1029:774], main_dev_inR1[773:262], main_dev_inR1[261:6], main_dev_inR1[5:0], main_dev_outR1);
  assign {__continue, __out0, __resumption_tag_next, __st0_next, __st1_next, __st2_next, __st3_next} = (zll_pure_dispatch6_in[1037:1036] == 2'h1) ? ((zll_main_loop125_in[5:0] == 6'h3f) ? main_dev_outR1 : main_loop_out) : ((zll_pure_dispatch8_in[1037:1036] == 2'h2) ? main_dev_out : ((zll_pure_dispatch16_in[1037:1036] == 2'h3) ? zll_main_dev89_outR1 : zll_main_dev89_out));
  initial {__resumption_tag, __st0, __st1, __st2, __st3} <= {1'h1, {11'h40d{1'h0}}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      {__resumption_tag, __st0, __st1, __st2, __st3} <= {1'h1, {11'h40d{1'h0}}};
    end else begin
      {__resumption_tag, __st0, __st1, __st2, __st3} <= {__resumption_tag_next, __st0_next, __st1_next, __st2_next, __st3_next};
    end
  end
endmodule

module ZLL_Main_dev89 (input logic [513:0] arg0,
  input logic [255:0] arg1,
  input logic [511:0] arg2,
  input logic [255:0] arg3,
  input logic [5:0] arg4,
  output logic [1296:0] res);
  logic [1029:0] main_loop_in;
  logic [1296:0] main_loop_out;
  assign main_loop_in = {arg1, arg2, arg3, arg4};
  Main_loop  inst (main_loop_in[1029:774], main_loop_in[773:262], main_loop_in[261:6], main_loop_in[5:0], main_loop_out);
  assign res = main_loop_out;
endmodule

module ZLL_Main_dev78 (input logic [511:0] arg0,
  input logic [255:0] arg1,
  input logic [511:0] arg2,
  input logic [255:0] arg3,
  input logic [5:0] arg4,
  output logic [1029:0] res);
  assign res = {arg1, arg0, arg3, arg4};
endmodule

module Main_dev (input logic [513:0] arg0,
  input logic [255:0] arg1,
  input logic [511:0] arg2,
  input logic [255:0] arg3,
  input logic [5:0] arg4,
  output logic [1296:0] res);
  logic [1543:0] zll_main_dev90_in;
  logic [1029:0] zll_main_dev63_in;
  logic [1285:0] zll_main_dev57_in;
  logic [1285:0] zll_main_dev65_in;
  logic [1285:0] zll_main_dev87_in;
  logic [1285:0] zll_main_dev10_in;
  logic [1285:0] zll_main_dev34_in;
  logic [1296:0] zll_main_dev91_in;
  logic [1296:0] zll_main_dev62_in;
  logic [1285:0] zll_main_dev12_in;
  logic [1285:0] zll_main_dev1_in;
  logic [1285:0] zll_main_dev9_in;
  logic [1543:0] zll_main_dev82_in;
  logic [1541:0] zll_main_dev44_in;
  logic [1541:0] zll_main_dev30_in;
  logic [1797:0] zll_main_dev38_in;
  logic [1797:0] zll_main_dev27_in;
  logic [1797:0] zll_main_dev41_in;
  logic [1797:0] zll_main_dev24_in;
  logic [1797:0] zll_main_dev49_in;
  logic [1797:0] zll_main_dev39_in;
  logic [1541:0] zll_main_dev20_in;
  logic [1541:0] zll_main_dev4_in;
  logic [1541:0] zll_main_dev52_in;
  logic [1541:0] zll_main_dev16_in;
  logic [1541:0] zll_main_dev51_in;
  logic [1541:0] zll_main_dev66_in;
  logic [1541:0] zll_main_dev22_in;
  logic [1541:0] zll_main_dev78_in;
  logic [1029:0] zll_main_dev78_out;
  logic [1029:0] zll_main_dev32_in;
  logic [1296:0] zll_main_dev32_out;
  logic [1296:0] zll_main_dev21_in;
  logic [1296:0] zll_main_dev80_in;
  logic [1029:0] zll_main_dev70_in;
  logic [1543:0] zll_main_dev74_in;
  logic [1541:0] zll_main_dev2_in;
  logic [1541:0] zll_main_dev25_in;
  logic [1541:0] zll_main_dev84_in;
  logic [1541:0] zll_main_dev59_in;
  logic [1541:0] zll_main_dev64_in;
  logic [1541:0] zll_main_dev92_in;
  logic [1541:0] zll_main_dev28_in;
  logic [1541:0] zll_main_dev61_in;
  logic [1797:0] zll_main_dev67_in;
  logic [1797:0] zll_main_dev6_in;
  logic [1797:0] zll_main_dev45_in;
  logic [1797:0] zll_main_dev75_in;
  logic [1797:0] zll_main_dev77_in;
  logic [1541:0] zll_main_dev14_in;
  logic [1541:0] zll_main_dev78_inR1;
  logic [1029:0] zll_main_dev78_outR1;
  logic [1029:0] zll_main_dev32_inR1;
  logic [1296:0] zll_main_dev32_outR1;
  logic [1296:0] zll_main_dev18_in;
  logic [1296:0] zll_main_dev13_in;
  logic [1029:0] zll_main_dev85_in;
  logic [1029:0] zll_main_dev72_in;
  logic [1029:0] zll_main_dev56_in;
  assign zll_main_dev90_in = {arg4, arg3, arg2, arg1, arg0};
  assign zll_main_dev63_in = {zll_main_dev90_in[769:514], zll_main_dev90_in[1281:770], zll_main_dev90_in[1537:1282], zll_main_dev90_in[1543:1538]};
  assign zll_main_dev57_in = {zll_main_dev63_in[261:6], zll_main_dev63_in[1029:774], zll_main_dev63_in[773:262], zll_main_dev63_in[261:6], zll_main_dev63_in[5:0]};
  assign zll_main_dev65_in = zll_main_dev57_in[1285:0];
  assign zll_main_dev87_in = {zll_main_dev65_in[1029:774], zll_main_dev65_in[1285:1030], zll_main_dev65_in[773:262], zll_main_dev65_in[261:6], zll_main_dev65_in[5:0]};
  assign zll_main_dev10_in = {zll_main_dev87_in[1285:1030], zll_main_dev87_in[773:262], zll_main_dev87_in[1029:774], zll_main_dev87_in[261:6], zll_main_dev87_in[5:0]};
  assign zll_main_dev34_in = {zll_main_dev10_in[1285:1030], zll_main_dev10_in[261:6], zll_main_dev10_in[1029:518], zll_main_dev10_in[517:262], zll_main_dev10_in[5:0]};
  assign zll_main_dev91_in = {11'h0, zll_main_dev34_in[261:6], zll_main_dev34_in[1285:1030], zll_main_dev34_in[773:262], zll_main_dev34_in[1029:774], zll_main_dev34_in[5:0]};
  assign zll_main_dev62_in = zll_main_dev91_in[1296:0];
  assign zll_main_dev12_in = {zll_main_dev62_in[1285:1030], zll_main_dev62_in[1029:774], zll_main_dev62_in[773:262], zll_main_dev62_in[261:6], zll_main_dev62_in[5:0]};
  assign zll_main_dev1_in = {zll_main_dev12_in[773:262], zll_main_dev12_in[1285:1030], zll_main_dev12_in[1029:774], zll_main_dev12_in[261:6], zll_main_dev12_in[5:0]};
  assign zll_main_dev9_in = {zll_main_dev1_in[773:518], zll_main_dev1_in[517:262], zll_main_dev1_in[1285:774], zll_main_dev1_in[261:6], zll_main_dev1_in[5:0]};
  assign zll_main_dev82_in = {arg4, arg3, arg2, arg1, arg0};
  assign zll_main_dev44_in = {zll_main_dev82_in[1543:1538], zll_main_dev82_in[1537:1282], zll_main_dev82_in[1281:770], zll_main_dev82_in[769:514], zll_main_dev82_in[511:0]};
  assign zll_main_dev30_in = {zll_main_dev44_in[511:0], zll_main_dev44_in[767:512], zll_main_dev44_in[1279:768], zll_main_dev44_in[1535:1280], zll_main_dev44_in[1541:1536]};
  assign zll_main_dev38_in = {zll_main_dev30_in[1541:1030], zll_main_dev30_in[261:6], zll_main_dev30_in[1029:774], zll_main_dev30_in[773:262], zll_main_dev30_in[261:6], zll_main_dev30_in[5:0]};
  assign zll_main_dev27_in = {zll_main_dev38_in[1797:1286], zll_main_dev38_in[1285:0]};
  assign zll_main_dev41_in = {zll_main_dev27_in[1285:1030], zll_main_dev27_in[1797:1286], zll_main_dev27_in[1029:774], zll_main_dev27_in[773:262], zll_main_dev27_in[261:6], zll_main_dev27_in[5:0]};
  assign zll_main_dev24_in = {zll_main_dev41_in[1029:774], zll_main_dev41_in[1797:1542], zll_main_dev41_in[1541:1030], zll_main_dev41_in[773:262], zll_main_dev41_in[261:6], zll_main_dev41_in[5:0]};
  assign zll_main_dev49_in = {zll_main_dev24_in[1797:1542], zll_main_dev24_in[1541:1286], zll_main_dev24_in[773:262], zll_main_dev24_in[1285:774], zll_main_dev24_in[261:6], zll_main_dev24_in[5:0]};
  assign zll_main_dev39_in = {zll_main_dev49_in[773:262], zll_main_dev49_in[1541:1286], zll_main_dev49_in[1797:1542], zll_main_dev49_in[1285:774], zll_main_dev49_in[261:6], zll_main_dev49_in[5:0]};
  assign zll_main_dev20_in = {zll_main_dev39_in[1797:1286], zll_main_dev39_in[1285:1030], zll_main_dev39_in[773:262], zll_main_dev39_in[261:6], zll_main_dev39_in[5:0]};
  assign zll_main_dev4_in = {zll_main_dev20_in[1541:1030], zll_main_dev20_in[1029:0]};
  assign zll_main_dev52_in = {zll_main_dev4_in[773:262], zll_main_dev4_in[1541:1030], zll_main_dev4_in[1029:774], zll_main_dev4_in[261:6], zll_main_dev4_in[5:0]};
  assign zll_main_dev16_in = {zll_main_dev52_in[1029:518], zll_main_dev52_in[517:262], zll_main_dev52_in[1541:1030], zll_main_dev52_in[261:6], zll_main_dev52_in[5:0]};
  assign zll_main_dev51_in = {zll_main_dev16_in[1541:1030], zll_main_dev16_in[1029:774], zll_main_dev16_in[773:262], zll_main_dev16_in[261:6], 6'h0};
  assign zll_main_dev66_in = {zll_main_dev51_in[1541:1030], zll_main_dev51_in[1029:0]};
  assign zll_main_dev22_in = {zll_main_dev66_in[773:262], zll_main_dev66_in[1541:1030], zll_main_dev66_in[1029:774], zll_main_dev66_in[261:6], zll_main_dev66_in[5:0]};
  assign zll_main_dev78_in = {zll_main_dev22_in[1029:518], zll_main_dev22_in[517:262], zll_main_dev22_in[1541:1030], zll_main_dev22_in[261:6], zll_main_dev22_in[5:0]};
  ZLL_Main_dev78  inst (zll_main_dev78_in[1541:1030], zll_main_dev78_in[1029:774], zll_main_dev78_in[773:262], zll_main_dev78_in[261:6], zll_main_dev78_in[5:0], zll_main_dev78_out);
  assign zll_main_dev32_in = zll_main_dev78_out;
  ZLL_Main_dev32  instR1 (zll_main_dev32_in[1029:0], zll_main_dev32_out);
  assign zll_main_dev21_in = zll_main_dev32_out;
  assign zll_main_dev80_in = zll_main_dev21_in[1296:0];
  assign zll_main_dev70_in = {zll_main_dev80_in[1029:774], zll_main_dev80_in[773:262], zll_main_dev80_in[261:6], zll_main_dev80_in[5:0]};
  assign zll_main_dev74_in = {arg4, arg3, arg2, arg1, arg0};
  assign zll_main_dev2_in = {zll_main_dev74_in[1543:1538], zll_main_dev74_in[1537:1282], zll_main_dev74_in[1281:770], zll_main_dev74_in[769:514], zll_main_dev74_in[511:0]};
  assign zll_main_dev25_in = {zll_main_dev2_in[511:0], zll_main_dev2_in[767:512], zll_main_dev2_in[1279:768], zll_main_dev2_in[1535:1280], zll_main_dev2_in[1541:1536]};
  assign zll_main_dev84_in = {zll_main_dev25_in[1541:1030], zll_main_dev25_in[1029:774], zll_main_dev25_in[773:262], 256'h6a09e667bb67ae853c6ef372a54ff53a510e527f9b05688c1f83d9ab5be0cd19, zll_main_dev25_in[5:0]};
  assign zll_main_dev59_in = {zll_main_dev84_in[1541:1030], zll_main_dev84_in[1029:0]};
  assign zll_main_dev64_in = {zll_main_dev59_in[773:262], zll_main_dev59_in[1541:1030], zll_main_dev59_in[1029:774], zll_main_dev59_in[261:6], zll_main_dev59_in[5:0]};
  assign zll_main_dev92_in = {zll_main_dev64_in[1029:518], zll_main_dev64_in[517:262], zll_main_dev64_in[1541:1030], zll_main_dev64_in[261:6], zll_main_dev64_in[5:0]};
  assign zll_main_dev28_in = {zll_main_dev92_in[1541:1030], zll_main_dev92_in[1029:774], zll_main_dev92_in[773:262], zll_main_dev92_in[261:6], 6'h0};
  assign zll_main_dev61_in = {zll_main_dev28_in[1541:1030], zll_main_dev28_in[1029:0]};
  assign zll_main_dev67_in = {zll_main_dev61_in[1541:1030], zll_main_dev61_in[261:6], zll_main_dev61_in[1029:774], zll_main_dev61_in[773:262], zll_main_dev61_in[261:6], zll_main_dev61_in[5:0]};
  assign zll_main_dev6_in = {zll_main_dev67_in[1797:1286], zll_main_dev67_in[1285:0]};
  assign zll_main_dev45_in = {zll_main_dev6_in[1797:1286], zll_main_dev6_in[1029:774], zll_main_dev6_in[1285:1030], zll_main_dev6_in[773:262], zll_main_dev6_in[261:6], zll_main_dev6_in[5:0]};
  assign zll_main_dev75_in = {zll_main_dev45_in[773:262], zll_main_dev45_in[1797:1286], zll_main_dev45_in[1285:1030], zll_main_dev45_in[1029:774], zll_main_dev45_in[261:6], zll_main_dev45_in[5:0]};
  assign zll_main_dev77_in = {zll_main_dev75_in[1285:774], zll_main_dev75_in[517:262], zll_main_dev75_in[773:518], zll_main_dev75_in[1797:1286], zll_main_dev75_in[261:6], zll_main_dev75_in[5:0]};
  assign zll_main_dev14_in = {zll_main_dev77_in[1797:1286], zll_main_dev77_in[1285:1030], zll_main_dev77_in[773:262], zll_main_dev77_in[261:6], zll_main_dev77_in[5:0]};
  assign zll_main_dev78_inR1 = {zll_main_dev14_in[1541:1030], zll_main_dev14_in[1029:0]};
  ZLL_Main_dev78  instR2 (zll_main_dev78_inR1[1541:1030], zll_main_dev78_inR1[1029:774], zll_main_dev78_inR1[773:262], zll_main_dev78_inR1[261:6], zll_main_dev78_inR1[5:0], zll_main_dev78_outR1);
  assign zll_main_dev32_inR1 = zll_main_dev78_outR1;
  ZLL_Main_dev32  instR3 (zll_main_dev32_inR1[1029:0], zll_main_dev32_outR1);
  assign zll_main_dev18_in = zll_main_dev32_outR1;
  assign zll_main_dev13_in = zll_main_dev18_in[1296:0];
  assign zll_main_dev85_in = {zll_main_dev13_in[1029:774], zll_main_dev13_in[773:262], zll_main_dev13_in[261:6], zll_main_dev13_in[5:0]};
  assign zll_main_dev72_in = {zll_main_dev85_in[773:262], zll_main_dev85_in[1029:774], zll_main_dev85_in[261:6], zll_main_dev85_in[5:0]};
  assign zll_main_dev56_in = {zll_main_dev72_in[517:262], zll_main_dev72_in[1029:518], zll_main_dev72_in[261:6], zll_main_dev72_in[5:0]};
  assign res = (zll_main_dev74_in[513:512] == 2'h0) ? {{3'h5, {9'h108{1'h0}}}, zll_main_dev56_in[1029:774], zll_main_dev56_in[773:262], zll_main_dev56_in[261:6], zll_main_dev56_in[5:0]} : ((zll_main_dev82_in[513:512] == 2'h1) ? {267'h50000000000000000000000000000000000000000000000000000000000000000c0, zll_main_dev70_in[1029:774], zll_main_dev70_in[773:262], zll_main_dev70_in[261:6], zll_main_dev70_in[5:0]} : {3'h4, zll_main_dev9_in[1285:1030], 8'h80, zll_main_dev9_in[1029:774], zll_main_dev9_in[773:262], zll_main_dev9_in[261:6], zll_main_dev9_in[5:0]});
endmodule

module Main_loop (input logic [255:0] arg0,
  input logic [511:0] arg1,
  input logic [255:0] arg2,
  input logic [5:0] arg3,
  output logic [1296:0] res);
  logic [1035:0] zll_main_loop148_in;
  logic [1035:0] zll_main_loop80_in;
  logic [1035:0] zll_main_loop128_in;
  logic [1035:0] zll_main_loop42_in;
  logic [1541:0] zll_main_loop45_in;
  logic [1541:0] zll_main_loop140_in;
  logic [1541:0] zll_main_loop97_in;
  logic [1541:0] zll_main_loop39_in;
  logic [2053:0] zll_main_loop40_in;
  logic [2053:0] zll_main_loop66_in;
  logic [2053:0] zll_main_loop101_in;
  logic [2053:0] zll_main_loop63_in;
  logic [2053:0] zll_main_loop49_in;
  logic [2053:0] zll_main_loop160_in;
  logic [2053:0] zll_main_loop156_in;
  logic [2053:0] zll_main_loop1_in;
  logic [2053:0] zll_main_loop123_in;
  logic [2053:0] zll_main_loop126_in;
  logic [2053:0] zll_main_loop144_in;
  logic [2053:0] zll_main_loop71_in;
  logic [2053:0] zll_main_loop64_in;
  logic [2053:0] zll_main_loop92_in;
  logic [2053:0] zll_main_loop124_in;
  logic [2053:0] zll_main_loop51_in;
  logic [2053:0] zll_main_loop46_in;
  logic [2053:0] zll_main_loop116_in;
  logic [2021:0] zll_main_loop96_in;
  logic [1989:0] zll_main_loop_in;
  logic [1957:0] zll_main_loop38_in;
  logic [1925:0] zll_main_loop54_in;
  logic [1893:0] zll_main_loop157_in;
  logic [1861:0] zll_main_loop11_in;
  logic [1829:0] zll_main_loop132_in;
  logic [1797:0] zll_main_loop77_in;
  logic [1765:0] zll_main_loop136_in;
  logic [1733:0] zll_main_loop150_in;
  logic [1701:0] zll_main_loop75_in;
  logic [1669:0] zll_main_loop19_in;
  logic [1637:0] zll_main_loop146_in;
  logic [1605:0] zll_main_loop141_in;
  logic [511:0] main_updatesched_in;
  logic [511:0] zll_main_updatesched4_in;
  logic [511:0] zll_main_updatesched13_in;
  logic [511:0] zll_main_updatesched3_in;
  logic [511:0] zll_main_updatesched15_in;
  logic [511:0] zll_main_updatesched7_in;
  logic [511:0] zll_main_updatesched5_in;
  logic [511:0] zll_main_updatesched_in;
  logic [511:0] zll_main_updatesched1_in;
  logic [511:0] zll_main_updatesched6_in;
  logic [511:0] zll_main_updatesched8_in;
  logic [511:0] zll_main_updatesched12_in;
  logic [511:0] zll_main_updatesched14_in;
  logic [511:0] zll_main_updatesched2_in;
  logic [31:0] main_sigma1_in;
  logic [31:0] main_rotater17_in;
  logic [31:0] zll_main_rotater1729_in;
  logic [31:0] zll_main_rotater1710_in;
  logic [31:0] zll_main_rotater1727_in;
  logic [31:0] zll_main_rotater1724_in;
  logic [31:0] zll_main_rotater1730_in;
  logic [31:0] zll_main_rotater178_in;
  logic [31:0] zll_main_rotater177_in;
  logic [31:0] zll_main_rotater175_in;
  logic [31:0] zll_main_rotater1714_in;
  logic [31:0] zll_main_rotater1721_in;
  logic [31:0] zll_main_rotater1712_in;
  logic [31:0] zll_main_rotater171_in;
  logic [31:0] zll_main_rotater1711_in;
  logic [31:0] zll_main_rotater1723_in;
  logic [31:0] zll_main_rotater1717_in;
  logic [31:0] zll_main_rotater1715_in;
  logic [31:0] zll_main_rotater1716_in;
  logic [31:0] zll_main_rotater179_in;
  logic [31:0] zll_main_rotater173_in;
  logic [31:0] zll_main_rotater1726_in;
  logic [31:0] zll_main_rotater176_in;
  logic [31:0] zll_main_rotater1713_in;
  logic [31:0] zll_main_rotater1728_in;
  logic [31:0] zll_main_rotater17_in;
  logic [31:0] zll_main_rotater1719_in;
  logic [31:0] zll_main_rotater174_in;
  logic [31:0] main_rotater19_in;
  logic [31:0] zll_main_rotater1931_in;
  logic [31:0] zll_main_rotater1912_in;
  logic [31:0] zll_main_rotater198_in;
  logic [31:0] zll_main_rotater1911_in;
  logic [31:0] zll_main_rotater1929_in;
  logic [31:0] zll_main_rotater194_in;
  logic [31:0] zll_main_rotater1930_in;
  logic [31:0] zll_main_rotater1918_in;
  logic [31:0] zll_main_rotater1920_in;
  logic [31:0] zll_main_rotater196_in;
  logic [31:0] zll_main_rotater1924_in;
  logic [31:0] zll_main_rotater1923_in;
  logic [31:0] zll_main_rotater1916_in;
  logic [31:0] zll_main_rotater1919_in;
  logic [31:0] zll_main_rotater1917_in;
  logic [31:0] zll_main_rotater1926_in;
  logic [31:0] zll_main_rotater195_in;
  logic [31:0] zll_main_rotater1914_in;
  logic [31:0] zll_main_rotater193_in;
  logic [31:0] zll_main_rotater192_in;
  logic [31:0] zll_main_rotater197_in;
  logic [31:0] zll_main_rotater19_in;
  logic [31:0] zll_main_rotater199_in;
  logic [31:0] zll_main_rotater1928_in;
  logic [31:0] zll_main_rotater1910_in;
  logic [63:0] xorw32_in;
  logic [31:0] extres;
  logic [31:0] main_shiftr10_in;
  logic [31:0] zll_main_shiftr1028_in;
  logic [31:0] zll_main_shiftr109_in;
  logic [31:0] zll_main_shiftr105_in;
  logic [31:0] zll_main_shiftr10_in;
  logic [31:0] zll_main_shiftr1013_in;
  logic [31:0] zll_main_shiftr108_in;
  logic [31:0] zll_main_shiftr1011_in;
  logic [31:0] zll_main_shiftr1016_in;
  logic [31:0] zll_main_shiftr1021_in;
  logic [31:0] zll_main_shiftr1024_in;
  logic [31:0] zll_main_shiftr103_in;
  logic [31:0] zll_main_shiftr106_in;
  logic [31:0] zll_main_shiftr1017_in;
  logic [31:0] zll_main_shiftr1012_in;
  logic [31:0] zll_main_shiftr1022_in;
  logic [31:0] zll_main_shiftr1030_in;
  logic [31:0] zll_main_shiftr104_in;
  logic [31:0] zll_main_shiftr1018_in;
  logic [30:0] zll_main_shiftr1020_in;
  logic [29:0] zll_main_shiftr107_in;
  logic [28:0] zll_main_shiftr1027_in;
  logic [27:0] zll_main_shiftr1026_in;
  logic [26:0] zll_main_shiftr1014_in;
  logic [25:0] zll_main_shiftr1015_in;
  logic [24:0] zll_main_shiftr1023_in;
  logic [23:0] zll_main_shiftr1010_in;
  logic [22:0] zll_main_shiftr101_in;
  logic [63:0] xorw32_inR1;
  logic [31:0] extresR1;
  logic [63:0] plusw32_in;
  logic [31:0] extresR2;
  logic [31:0] main_sigma0_in;
  logic [31:0] main_rotater7_in;
  logic [31:0] zll_main_rotater713_in;
  logic [31:0] zll_main_rotater7_in;
  logic [31:0] zll_main_rotater727_in;
  logic [31:0] zll_main_rotater76_in;
  logic [31:0] zll_main_rotater722_in;
  logic [31:0] zll_main_rotater725_in;
  logic [31:0] zll_main_rotater71_in;
  logic [31:0] zll_main_rotater75_in;
  logic [31:0] zll_main_rotater719_in;
  logic [31:0] zll_main_rotater728_in;
  logic [31:0] zll_main_rotater717_in;
  logic [31:0] zll_main_rotater731_in;
  logic [31:0] zll_main_rotater724_in;
  logic [31:0] zll_main_rotater711_in;
  logic [31:0] zll_main_rotater72_in;
  logic [31:0] zll_main_rotater720_in;
  logic [31:0] zll_main_rotater718_in;
  logic [31:0] zll_main_rotater79_in;
  logic [31:0] zll_main_rotater714_in;
  logic [31:0] zll_main_rotater74_in;
  logic [31:0] zll_main_rotater77_in;
  logic [31:0] zll_main_rotater712_in;
  logic [31:0] zll_main_rotater721_in;
  logic [31:0] zll_main_rotater729_in;
  logic [31:0] zll_main_rotater726_in;
  logic [31:0] zll_main_rotater73_in;
  logic [31:0] zll_main_rotater78_in;
  logic [31:0] zll_main_rotater716_in;
  logic [31:0] zll_main_rotater715_in;
  logic [31:0] main_rotater18_in;
  logic [31:0] zll_main_rotater1825_in;
  logic [31:0] zll_main_rotater1818_in;
  logic [31:0] zll_main_rotater1828_in;
  logic [31:0] zll_main_rotater1826_in;
  logic [31:0] zll_main_rotater1824_in;
  logic [31:0] zll_main_rotater188_in;
  logic [31:0] zll_main_rotater1817_in;
  logic [31:0] zll_main_rotater181_in;
  logic [31:0] zll_main_rotater1811_in;
  logic [31:0] zll_main_rotater1830_in;
  logic [31:0] zll_main_rotater1821_in;
  logic [31:0] zll_main_rotater1813_in;
  logic [31:0] zll_main_rotater186_in;
  logic [31:0] zll_main_rotater1827_in;
  logic [31:0] zll_main_rotater185_in;
  logic [31:0] zll_main_rotater1820_in;
  logic [31:0] zll_main_rotater1822_in;
  logic [31:0] zll_main_rotater1814_in;
  logic [31:0] zll_main_rotater1815_in;
  logic [31:0] zll_main_rotater184_in;
  logic [31:0] zll_main_rotater182_in;
  logic [31:0] zll_main_rotater1823_in;
  logic [31:0] zll_main_rotater1829_in;
  logic [31:0] zll_main_rotater1810_in;
  logic [31:0] zll_main_rotater183_in;
  logic [31:0] zll_main_rotater1816_in;
  logic [31:0] zll_main_rotater189_in;
  logic [31:0] zll_main_rotater18_in;
  logic [31:0] zll_main_rotater1812_in;
  logic [63:0] xorw32_inR2;
  logic [31:0] extresR3;
  logic [31:0] main_shiftr3_in;
  logic [31:0] zll_main_shiftr311_in;
  logic [31:0] zll_main_shiftr38_in;
  logic [31:0] zll_main_shiftr330_in;
  logic [31:0] zll_main_shiftr36_in;
  logic [31:0] zll_main_shiftr312_in;
  logic [31:0] zll_main_shiftr326_in;
  logic [31:0] zll_main_shiftr322_in;
  logic [31:0] zll_main_shiftr321_in;
  logic [31:0] zll_main_shiftr316_in;
  logic [31:0] zll_main_shiftr323_in;
  logic [31:0] zll_main_shiftr3_in;
  logic [31:0] zll_main_shiftr33_in;
  logic [31:0] zll_main_shiftr310_in;
  logic [31:0] zll_main_shiftr39_in;
  logic [31:0] zll_main_shiftr320_in;
  logic [31:0] zll_main_shiftr327_in;
  logic [31:0] zll_main_shiftr315_in;
  logic [31:0] zll_main_shiftr329_in;
  logic [31:0] zll_main_shiftr331_in;
  logic [31:0] zll_main_shiftr324_in;
  logic [31:0] zll_main_shiftr32_in;
  logic [31:0] zll_main_shiftr325_in;
  logic [31:0] zll_main_shiftr314_in;
  logic [31:0] zll_main_shiftr35_in;
  logic [31:0] zll_main_shiftr31_in;
  logic [31:0] zll_main_shiftr37_in;
  logic [31:0] zll_main_shiftr313_in;
  logic [30:0] zll_main_shiftr328_in;
  logic [29:0] zll_main_shiftr34_in;
  logic [63:0] xorw32_inR3;
  logic [31:0] extresR4;
  logic [63:0] plusw32_inR1;
  logic [31:0] extresR5;
  logic [63:0] plusw32_inR2;
  logic [31:0] extresR6;
  logic [1061:0] zll_main_loop74_in;
  logic [1061:0] zll_main_loop58_in;
  logic [1061:0] zll_main_loop17_in;
  logic [1067:0] zll_main_loop151_in;
  logic [1067:0] zll_main_loop20_in;
  logic [1067:0] zll_main_loop32_in;
  logic [1067:0] zll_main_loop103_in;
  logic [1067:0] zll_main_loop72_in;
  logic [1323:0] zll_main_loop15_in;
  logic [1323:0] zll_main_loop60_in;
  logic [1323:0] zll_main_loop3_in;
  logic [1323:0] zll_main_loop5_in;
  logic [1323:0] zll_main_loop35_in;
  logic [5:0] main_seed_in;
  logic [5:0] lit_in;
  logic [5:0] lit_inR1;
  logic [5:0] lit_inR2;
  logic [5:0] lit_inR3;
  logic [5:0] lit_inR4;
  logic [5:0] lit_inR5;
  logic [5:0] lit_inR6;
  logic [5:0] lit_inR7;
  logic [5:0] lit_inR8;
  logic [5:0] lit_inR9;
  logic [5:0] lit_inR10;
  logic [5:0] lit_inR11;
  logic [5:0] lit_inR12;
  logic [5:0] lit_inR13;
  logic [5:0] lit_inR14;
  logic [5:0] lit_inR15;
  logic [5:0] lit_inR16;
  logic [5:0] lit_inR17;
  logic [5:0] lit_inR18;
  logic [5:0] lit_inR19;
  logic [5:0] lit_inR20;
  logic [5:0] lit_inR21;
  logic [5:0] lit_inR22;
  logic [5:0] lit_inR23;
  logic [5:0] lit_inR24;
  logic [5:0] lit_inR25;
  logic [5:0] lit_inR26;
  logic [5:0] lit_inR27;
  logic [5:0] lit_inR28;
  logic [5:0] lit_inR29;
  logic [5:0] lit_inR30;
  logic [5:0] lit_inR31;
  logic [5:0] lit_inR32;
  logic [5:0] lit_inR33;
  logic [5:0] lit_inR34;
  logic [5:0] lit_inR35;
  logic [5:0] lit_inR36;
  logic [5:0] lit_inR37;
  logic [5:0] lit_inR38;
  logic [5:0] lit_inR39;
  logic [5:0] lit_inR40;
  logic [5:0] lit_inR41;
  logic [5:0] lit_inR42;
  logic [5:0] lit_inR43;
  logic [5:0] lit_inR44;
  logic [5:0] lit_inR45;
  logic [5:0] lit_inR46;
  logic [5:0] lit_inR47;
  logic [5:0] lit_inR48;
  logic [5:0] lit_inR49;
  logic [5:0] lit_inR50;
  logic [5:0] lit_inR51;
  logic [5:0] lit_inR52;
  logic [5:0] lit_inR53;
  logic [5:0] lit_inR54;
  logic [5:0] lit_inR55;
  logic [5:0] lit_inR56;
  logic [5:0] lit_inR57;
  logic [5:0] lit_inR58;
  logic [5:0] lit_inR59;
  logic [5:0] lit_inR60;
  logic [5:0] lit_inR61;
  logic [5:0] lit_inR62;
  logic [319:0] main_step256_in;
  logic [319:0] zll_main_step2568_in;
  logic [319:0] zll_main_step2562_in;
  logic [319:0] zll_main_step2561_in;
  logic [319:0] zll_main_step256_in;
  logic [319:0] zll_main_step2565_in;
  logic [319:0] zll_main_step2566_in;
  logic [31:0] main_bigsigma1_in;
  logic [31:0] main_bigsigma1_out;
  logic [95:0] main_ch_in;
  logic [31:0] main_ch_out;
  logic [63:0] plusw32_inR3;
  logic [31:0] extresR7;
  logic [63:0] plusw32_inR4;
  logic [31:0] extresR8;
  logic [63:0] plusw32_inR5;
  logic [31:0] extresR9;
  logic [63:0] plusw32_inR6;
  logic [31:0] extresR10;
  logic [31:0] main_bigsigma0_in;
  logic [31:0] main_rotater2_in;
  logic [31:0] zll_main_rotater211_in;
  logic [31:0] zll_main_rotater210_in;
  logic [31:0] zll_main_rotater213_in;
  logic [31:0] zll_main_rotater23_in;
  logic [31:0] zll_main_rotater242_in;
  logic [31:0] zll_main_rotater220_in;
  logic [31:0] zll_main_rotater24_in;
  logic [31:0] zll_main_rotater233_in;
  logic [31:0] zll_main_rotater212_in;
  logic [31:0] zll_main_rotater235_in;
  logic [31:0] zll_main_rotater230_in;
  logic [31:0] zll_main_rotater26_in;
  logic [31:0] zll_main_rotater232_in;
  logic [31:0] zll_main_rotater236_in;
  logic [31:0] zll_main_rotater216_in;
  logic [31:0] zll_main_rotater241_in;
  logic [31:0] zll_main_rotater29_in;
  logic [31:0] zll_main_rotater218_in;
  logic [31:0] zll_main_rotater239_in;
  logic [31:0] zll_main_rotater231_in;
  logic [31:0] zll_main_rotater28_in;
  logic [31:0] zll_main_rotater215_in;
  logic [31:0] zll_main_rotater219_in;
  logic [31:0] zll_main_rotater27_in;
  logic [31:0] zll_main_rotater214_in;
  logic [31:0] zll_main_rotater217_in;
  logic [31:0] zll_main_rotater240_in;
  logic [31:0] zll_main_rotater2_in;
  logic [31:0] zll_main_rotater237_in;
  logic [31:0] main_rotater13_in;
  logic [31:0] zll_main_rotater1323_in;
  logic [31:0] zll_main_rotater1316_in;
  logic [31:0] zll_main_rotater1328_in;
  logic [31:0] zll_main_rotater1317_in;
  logic [31:0] zll_main_rotater1321_in;
  logic [31:0] zll_main_rotater1319_in;
  logic [31:0] zll_main_rotater1326_in;
  logic [31:0] zll_main_rotater1331_in;
  logic [31:0] zll_main_rotater1310_in;
  logic [31:0] zll_main_rotater1311_in;
  logic [31:0] zll_main_rotater131_in;
  logic [31:0] zll_main_rotater1325_in;
  logic [31:0] zll_main_rotater1329_in;
  logic [31:0] zll_main_rotater1312_in;
  logic [31:0] zll_main_rotater132_in;
  logic [31:0] zll_main_rotater1327_in;
  logic [31:0] zll_main_rotater1322_in;
  logic [31:0] zll_main_rotater137_in;
  logic [31:0] zll_main_rotater134_in;
  logic [31:0] zll_main_rotater1330_in;
  logic [31:0] zll_main_rotater1320_in;
  logic [31:0] zll_main_rotater1315_in;
  logic [31:0] zll_main_rotater1313_in;
  logic [31:0] zll_main_rotater13_in;
  logic [31:0] zll_main_rotater136_in;
  logic [31:0] zll_main_rotater1318_in;
  logic [31:0] zll_main_rotater135_in;
  logic [31:0] zll_main_rotater133_in;
  logic [31:0] zll_main_rotater1314_in;
  logic [63:0] xorw32_inR4;
  logic [31:0] extresR11;
  logic [31:0] main_rotater22_in;
  logic [31:0] zll_main_rotater227_in;
  logic [31:0] zll_main_rotater2213_in;
  logic [31:0] zll_main_rotater2229_in;
  logic [31:0] zll_main_rotater2230_in;
  logic [31:0] zll_main_rotater2214_in;
  logic [31:0] zll_main_rotater2226_in;
  logic [31:0] zll_main_rotater2228_in;
  logic [31:0] zll_main_rotater221_in;
  logic [31:0] zll_main_rotater2224_in;
  logic [31:0] zll_main_rotater2211_in;
  logic [31:0] zll_main_rotater224_in;
  logic [31:0] zll_main_rotater2219_in;
  logic [31:0] zll_main_rotater2222_in;
  logic [31:0] zll_main_rotater229_in;
  logic [31:0] zll_main_rotater228_in;
  logic [31:0] zll_main_rotater22_in;
  logic [31:0] zll_main_rotater223_in;
  logic [31:0] zll_main_rotater2212_in;
  logic [31:0] zll_main_rotater2231_in;
  logic [31:0] zll_main_rotater222_in;
  logic [31:0] zll_main_rotater2227_in;
  logic [31:0] zll_main_rotater2210_in;
  logic [31:0] zll_main_rotater225_in;
  logic [31:0] zll_main_rotater226_in;
  logic [31:0] zll_main_rotater2216_in;
  logic [31:0] zll_main_rotater2220_in;
  logic [31:0] zll_main_rotater2217_in;
  logic [31:0] zll_main_rotater2221_in;
  logic [63:0] xorw32_inR5;
  logic [31:0] extresR12;
  logic [95:0] main_maj_in;
  logic [63:0] andw32_in;
  logic [31:0] extresR13;
  logic [63:0] andw32_inR1;
  logic [31:0] extresR14;
  logic [63:0] xorw32_inR6;
  logic [31:0] extresR15;
  logic [63:0] andw32_inR2;
  logic [31:0] extresR16;
  logic [63:0] xorw32_inR7;
  logic [31:0] extresR17;
  logic [63:0] plusw32_inR7;
  logic [31:0] extresR18;
  logic [63:0] plusw32_inR8;
  logic [31:0] extresR19;
  logic [31:0] main_bigsigma1_inR1;
  logic [31:0] main_bigsigma1_outR1;
  logic [95:0] main_ch_inR1;
  logic [31:0] main_ch_outR1;
  logic [63:0] plusw32_inR9;
  logic [31:0] extresR20;
  logic [63:0] plusw32_inR10;
  logic [31:0] extresR21;
  logic [63:0] plusw32_inR11;
  logic [31:0] extresR22;
  logic [63:0] plusw32_inR12;
  logic [31:0] extresR23;
  logic [63:0] plusw32_inR13;
  logic [31:0] extresR24;
  logic [1035:0] zll_main_loop6_in;
  logic [1035:0] zll_main_loop109_in;
  logic [1035:0] zll_main_loop107_in;
  logic [1035:0] zll_main_loop84_in;
  logic [5:0] main_incctr_in;
  logic [5:0] lit_inR63;
  logic [5:0] lit_inR64;
  logic [5:0] lit_inR65;
  logic [5:0] lit_inR66;
  logic [5:0] lit_inR67;
  logic [5:0] lit_inR68;
  logic [5:0] lit_inR69;
  logic [5:0] lit_inR70;
  logic [5:0] lit_inR71;
  logic [5:0] lit_inR72;
  logic [5:0] lit_inR73;
  logic [5:0] lit_inR74;
  logic [5:0] lit_inR75;
  logic [5:0] lit_inR76;
  logic [5:0] lit_inR77;
  logic [5:0] lit_inR78;
  logic [5:0] lit_inR79;
  logic [5:0] lit_inR80;
  logic [5:0] lit_inR81;
  logic [5:0] lit_inR82;
  logic [5:0] lit_inR83;
  logic [5:0] lit_inR84;
  logic [5:0] lit_inR85;
  logic [5:0] lit_inR86;
  logic [5:0] lit_inR87;
  logic [5:0] lit_inR88;
  logic [5:0] lit_inR89;
  logic [5:0] lit_inR90;
  logic [5:0] lit_inR91;
  logic [5:0] lit_inR92;
  logic [5:0] lit_inR93;
  logic [5:0] lit_inR94;
  logic [5:0] lit_inR95;
  logic [5:0] lit_inR96;
  logic [5:0] lit_inR97;
  logic [5:0] lit_inR98;
  logic [5:0] lit_inR99;
  logic [5:0] lit_inR100;
  logic [5:0] lit_inR101;
  logic [5:0] lit_inR102;
  logic [5:0] lit_inR103;
  logic [5:0] lit_inR104;
  logic [5:0] lit_inR105;
  logic [5:0] lit_inR106;
  logic [5:0] lit_inR107;
  logic [5:0] lit_inR108;
  logic [5:0] lit_inR109;
  logic [5:0] lit_inR110;
  logic [5:0] lit_inR111;
  logic [5:0] lit_inR112;
  logic [5:0] lit_inR113;
  logic [5:0] lit_inR114;
  logic [5:0] lit_inR115;
  logic [5:0] lit_inR116;
  logic [5:0] lit_inR117;
  logic [5:0] lit_inR118;
  logic [5:0] lit_inR119;
  logic [5:0] lit_inR120;
  logic [5:0] lit_inR121;
  logic [5:0] lit_inR122;
  logic [5:0] lit_inR123;
  logic [5:0] lit_inR124;
  logic [5:0] lit_inR125;
  logic [1035:0] zll_main_loop108_in;
  logic [1035:0] zll_main_loop8_in;
  logic [1035:0] zll_main_loop67_in;
  logic [1035:0] zll_main_loop55_in;
  logic [1035:0] zll_main_loop29_in;
  logic [1035:0] zll_main_loop112_in;
  logic [1035:0] zll_main_loop18_in;
  logic [1035:0] zll_main_loop122_in;
  logic [1296:0] zll_main_loop41_in;
  logic [1296:0] zll_main_loop162_in;
  logic [1035:0] zll_main_loop154_in;
  logic [1035:0] zll_main_loop111_in;
  logic [1035:0] zll_main_loop79_in;
  assign zll_main_loop148_in = {arg3, arg0, arg1, arg2, arg3};
  assign zll_main_loop80_in = zll_main_loop148_in[1035:0];
  assign zll_main_loop128_in = {zll_main_loop80_in[1035:1030], zll_main_loop80_in[773:262], zll_main_loop80_in[1029:774], zll_main_loop80_in[261:6], zll_main_loop80_in[5:0]};
  assign zll_main_loop42_in = {zll_main_loop128_in[1035:1030], zll_main_loop128_in[517:262], zll_main_loop128_in[1029:518], zll_main_loop128_in[261:6], zll_main_loop128_in[5:0]};
  assign zll_main_loop45_in = {zll_main_loop42_in[773:262], zll_main_loop42_in[1029:774], zll_main_loop42_in[773:262], zll_main_loop42_in[261:6], zll_main_loop42_in[5:0]};
  assign zll_main_loop140_in = zll_main_loop45_in[1541:0];
  assign zll_main_loop97_in = {zll_main_loop140_in[1029:774], zll_main_loop140_in[1541:1030], zll_main_loop140_in[773:262], zll_main_loop140_in[261:6], zll_main_loop140_in[5:0]};
  assign zll_main_loop39_in = {zll_main_loop97_in[1285:774], zll_main_loop97_in[1541:1286], zll_main_loop97_in[773:262], zll_main_loop97_in[261:6], zll_main_loop97_in[5:0]};
  assign zll_main_loop40_in = {zll_main_loop39_in[1029:774], zll_main_loop39_in[773:262], zll_main_loop39_in[5:0], zll_main_loop39_in[261:6], zll_main_loop39_in[1541:1030], zll_main_loop39_in[1541:1030]};
  assign zll_main_loop66_in = {zll_main_loop40_in[2053:1798], zll_main_loop40_in[1023:512], zll_main_loop40_in[1797:1286], zll_main_loop40_in[1285:1280], zll_main_loop40_in[1279:1024], zll_main_loop40_in[511:480], zll_main_loop40_in[479:448], zll_main_loop40_in[447:416], zll_main_loop40_in[415:384], zll_main_loop40_in[383:352], zll_main_loop40_in[351:320], zll_main_loop40_in[319:288], zll_main_loop40_in[287:256], zll_main_loop40_in[255:224], zll_main_loop40_in[223:192], zll_main_loop40_in[191:160], zll_main_loop40_in[159:128], zll_main_loop40_in[127:96], zll_main_loop40_in[95:64], zll_main_loop40_in[63:32], zll_main_loop40_in[31:0]};
  assign zll_main_loop101_in = {zll_main_loop66_in[2053:1798], zll_main_loop66_in[1797:1286], zll_main_loop66_in[1285:774], zll_main_loop66_in[511:480], zll_main_loop66_in[773:768], zll_main_loop66_in[767:512], zll_main_loop66_in[479:448], zll_main_loop66_in[447:416], zll_main_loop66_in[415:384], zll_main_loop66_in[383:352], zll_main_loop66_in[351:320], zll_main_loop66_in[319:288], zll_main_loop66_in[287:256], zll_main_loop66_in[255:224], zll_main_loop66_in[223:192], zll_main_loop66_in[191:160], zll_main_loop66_in[159:128], zll_main_loop66_in[127:96], zll_main_loop66_in[95:64], zll_main_loop66_in[63:32], zll_main_loop66_in[31:0]};
  assign zll_main_loop63_in = {zll_main_loop101_in[2053:1798], zll_main_loop101_in[1797:1286], zll_main_loop101_in[1285:774], zll_main_loop101_in[773:742], zll_main_loop101_in[741:736], zll_main_loop101_in[479:448], zll_main_loop101_in[735:480], zll_main_loop101_in[447:416], zll_main_loop101_in[415:384], zll_main_loop101_in[383:352], zll_main_loop101_in[351:320], zll_main_loop101_in[319:288], zll_main_loop101_in[287:256], zll_main_loop101_in[255:224], zll_main_loop101_in[223:192], zll_main_loop101_in[191:160], zll_main_loop101_in[159:128], zll_main_loop101_in[127:96], zll_main_loop101_in[95:64], zll_main_loop101_in[63:32], zll_main_loop101_in[31:0]};
  assign zll_main_loop49_in = {zll_main_loop63_in[2053:1798], zll_main_loop63_in[1797:1286], zll_main_loop63_in[1285:774], zll_main_loop63_in[773:742], zll_main_loop63_in[741:736], zll_main_loop63_in[447:416], zll_main_loop63_in[735:704], zll_main_loop63_in[703:448], zll_main_loop63_in[415:384], zll_main_loop63_in[383:352], zll_main_loop63_in[351:320], zll_main_loop63_in[319:288], zll_main_loop63_in[287:256], zll_main_loop63_in[255:224], zll_main_loop63_in[223:192], zll_main_loop63_in[191:160], zll_main_loop63_in[159:128], zll_main_loop63_in[127:96], zll_main_loop63_in[95:64], zll_main_loop63_in[63:32], zll_main_loop63_in[31:0]};
  assign zll_main_loop160_in = {zll_main_loop49_in[2053:1798], zll_main_loop49_in[1797:1286], zll_main_loop49_in[415:384], zll_main_loop49_in[1285:774], zll_main_loop49_in[773:742], zll_main_loop49_in[741:736], zll_main_loop49_in[735:704], zll_main_loop49_in[703:672], zll_main_loop49_in[671:416], zll_main_loop49_in[383:352], zll_main_loop49_in[351:320], zll_main_loop49_in[319:288], zll_main_loop49_in[287:256], zll_main_loop49_in[255:224], zll_main_loop49_in[223:192], zll_main_loop49_in[191:160], zll_main_loop49_in[159:128], zll_main_loop49_in[127:96], zll_main_loop49_in[95:64], zll_main_loop49_in[63:32], zll_main_loop49_in[31:0]};
  assign zll_main_loop156_in = {zll_main_loop160_in[2053:1798], zll_main_loop160_in[1797:1286], zll_main_loop160_in[1285:1254], zll_main_loop160_in[1253:742], zll_main_loop160_in[383:352], zll_main_loop160_in[741:710], zll_main_loop160_in[709:704], zll_main_loop160_in[703:672], zll_main_loop160_in[671:640], zll_main_loop160_in[639:384], zll_main_loop160_in[351:320], zll_main_loop160_in[319:288], zll_main_loop160_in[287:256], zll_main_loop160_in[255:224], zll_main_loop160_in[223:192], zll_main_loop160_in[191:160], zll_main_loop160_in[159:128], zll_main_loop160_in[127:96], zll_main_loop160_in[95:64], zll_main_loop160_in[63:32], zll_main_loop160_in[31:0]};
  assign zll_main_loop1_in = {zll_main_loop156_in[2053:1798], zll_main_loop156_in[351:320], zll_main_loop156_in[1797:1286], zll_main_loop156_in[1285:1254], zll_main_loop156_in[1253:742], zll_main_loop156_in[741:710], zll_main_loop156_in[709:678], zll_main_loop156_in[677:672], zll_main_loop156_in[671:640], zll_main_loop156_in[639:608], zll_main_loop156_in[607:352], zll_main_loop156_in[319:288], zll_main_loop156_in[287:256], zll_main_loop156_in[255:224], zll_main_loop156_in[223:192], zll_main_loop156_in[191:160], zll_main_loop156_in[159:128], zll_main_loop156_in[127:96], zll_main_loop156_in[95:64], zll_main_loop156_in[63:32], zll_main_loop156_in[31:0]};
  assign zll_main_loop123_in = {zll_main_loop1_in[2053:1798], zll_main_loop1_in[1797:1766], zll_main_loop1_in[1765:1254], zll_main_loop1_in[1253:1222], zll_main_loop1_in[1221:710], zll_main_loop1_in[709:678], zll_main_loop1_in[677:646], zll_main_loop1_in[645:640], zll_main_loop1_in[639:608], zll_main_loop1_in[607:576], zll_main_loop1_in[319:288], zll_main_loop1_in[575:320], zll_main_loop1_in[287:256], zll_main_loop1_in[255:224], zll_main_loop1_in[223:192], zll_main_loop1_in[191:160], zll_main_loop1_in[159:128], zll_main_loop1_in[127:96], zll_main_loop1_in[95:64], zll_main_loop1_in[63:32], zll_main_loop1_in[31:0]};
  assign zll_main_loop126_in = {zll_main_loop123_in[2053:1798], zll_main_loop123_in[1797:1766], zll_main_loop123_in[1765:1254], zll_main_loop123_in[1253:1222], zll_main_loop123_in[1221:710], zll_main_loop123_in[709:678], zll_main_loop123_in[287:256], zll_main_loop123_in[677:646], zll_main_loop123_in[645:640], zll_main_loop123_in[639:608], zll_main_loop123_in[607:576], zll_main_loop123_in[575:544], zll_main_loop123_in[543:288], zll_main_loop123_in[255:224], zll_main_loop123_in[223:192], zll_main_loop123_in[191:160], zll_main_loop123_in[159:128], zll_main_loop123_in[127:96], zll_main_loop123_in[95:64], zll_main_loop123_in[63:32], zll_main_loop123_in[31:0]};
  assign zll_main_loop144_in = {zll_main_loop126_in[2053:1798], zll_main_loop126_in[1797:1766], zll_main_loop126_in[1765:1254], zll_main_loop126_in[1253:1222], zll_main_loop126_in[1221:710], zll_main_loop126_in[709:678], zll_main_loop126_in[677:646], zll_main_loop126_in[645:614], zll_main_loop126_in[613:608], zll_main_loop126_in[255:224], zll_main_loop126_in[607:576], zll_main_loop126_in[575:544], zll_main_loop126_in[543:512], zll_main_loop126_in[511:256], zll_main_loop126_in[223:192], zll_main_loop126_in[191:160], zll_main_loop126_in[159:128], zll_main_loop126_in[127:96], zll_main_loop126_in[95:64], zll_main_loop126_in[63:32], zll_main_loop126_in[31:0]};
  assign zll_main_loop71_in = {zll_main_loop144_in[2053:1798], zll_main_loop144_in[1797:1766], zll_main_loop144_in[223:192], zll_main_loop144_in[1765:1254], zll_main_loop144_in[1253:1222], zll_main_loop144_in[1221:710], zll_main_loop144_in[709:678], zll_main_loop144_in[677:646], zll_main_loop144_in[645:614], zll_main_loop144_in[613:608], zll_main_loop144_in[607:576], zll_main_loop144_in[575:544], zll_main_loop144_in[543:512], zll_main_loop144_in[511:480], zll_main_loop144_in[479:224], zll_main_loop144_in[191:160], zll_main_loop144_in[159:128], zll_main_loop144_in[127:96], zll_main_loop144_in[95:64], zll_main_loop144_in[63:32], zll_main_loop144_in[31:0]};
  assign zll_main_loop64_in = {zll_main_loop71_in[2053:1798], zll_main_loop71_in[1797:1766], zll_main_loop71_in[1765:1734], zll_main_loop71_in[1733:1222], zll_main_loop71_in[1221:1190], zll_main_loop71_in[1189:678], zll_main_loop71_in[677:646], zll_main_loop71_in[645:614], zll_main_loop71_in[613:582], zll_main_loop71_in[191:160], zll_main_loop71_in[581:576], zll_main_loop71_in[575:544], zll_main_loop71_in[543:512], zll_main_loop71_in[511:480], zll_main_loop71_in[479:448], zll_main_loop71_in[447:192], zll_main_loop71_in[159:128], zll_main_loop71_in[127:96], zll_main_loop71_in[95:64], zll_main_loop71_in[63:32], zll_main_loop71_in[31:0]};
  assign zll_main_loop92_in = {zll_main_loop64_in[2053:1798], zll_main_loop64_in[1797:1766], zll_main_loop64_in[1765:1734], zll_main_loop64_in[1733:1222], zll_main_loop64_in[1221:1190], zll_main_loop64_in[1189:678], zll_main_loop64_in[159:128], zll_main_loop64_in[677:646], zll_main_loop64_in[645:614], zll_main_loop64_in[613:582], zll_main_loop64_in[581:550], zll_main_loop64_in[549:544], zll_main_loop64_in[543:512], zll_main_loop64_in[511:480], zll_main_loop64_in[479:448], zll_main_loop64_in[447:416], zll_main_loop64_in[415:160], zll_main_loop64_in[127:96], zll_main_loop64_in[95:64], zll_main_loop64_in[63:32], zll_main_loop64_in[31:0]};
  assign zll_main_loop124_in = {zll_main_loop92_in[2053:1798], zll_main_loop92_in[1797:1766], zll_main_loop92_in[1765:1734], zll_main_loop92_in[1733:1222], zll_main_loop92_in[1221:1190], zll_main_loop92_in[1189:678], zll_main_loop92_in[677:646], zll_main_loop92_in[645:614], zll_main_loop92_in[613:582], zll_main_loop92_in[581:550], zll_main_loop92_in[549:518], zll_main_loop92_in[517:512], zll_main_loop92_in[127:96], zll_main_loop92_in[511:480], zll_main_loop92_in[479:448], zll_main_loop92_in[447:416], zll_main_loop92_in[415:384], zll_main_loop92_in[383:128], zll_main_loop92_in[95:64], zll_main_loop92_in[63:32], zll_main_loop92_in[31:0]};
  assign zll_main_loop51_in = {zll_main_loop124_in[2053:1798], zll_main_loop124_in[1797:1766], zll_main_loop124_in[1765:1734], zll_main_loop124_in[1733:1222], zll_main_loop124_in[1221:1190], zll_main_loop124_in[1189:678], zll_main_loop124_in[677:646], zll_main_loop124_in[645:614], zll_main_loop124_in[613:582], zll_main_loop124_in[581:550], zll_main_loop124_in[549:518], zll_main_loop124_in[517:512], zll_main_loop124_in[511:480], zll_main_loop124_in[95:64], zll_main_loop124_in[479:448], zll_main_loop124_in[447:416], zll_main_loop124_in[415:384], zll_main_loop124_in[383:352], zll_main_loop124_in[351:96], zll_main_loop124_in[63:32], zll_main_loop124_in[31:0]};
  assign zll_main_loop46_in = {zll_main_loop51_in[2053:1798], zll_main_loop51_in[1797:1766], zll_main_loop51_in[1765:1734], zll_main_loop51_in[1733:1222], zll_main_loop51_in[1221:1190], zll_main_loop51_in[63:32], zll_main_loop51_in[1189:678], zll_main_loop51_in[677:646], zll_main_loop51_in[645:614], zll_main_loop51_in[613:582], zll_main_loop51_in[581:550], zll_main_loop51_in[549:518], zll_main_loop51_in[517:512], zll_main_loop51_in[511:480], zll_main_loop51_in[479:448], zll_main_loop51_in[447:416], zll_main_loop51_in[415:384], zll_main_loop51_in[383:352], zll_main_loop51_in[351:320], zll_main_loop51_in[319:64], zll_main_loop51_in[31:0]};
  assign zll_main_loop116_in = {zll_main_loop46_in[1733:1222], zll_main_loop46_in[549:518], zll_main_loop46_in[351:320], zll_main_loop46_in[383:352], zll_main_loop46_in[1221:1190], zll_main_loop46_in[613:582], zll_main_loop46_in[1797:1766], zll_main_loop46_in[319:288], zll_main_loop46_in[581:550], zll_main_loop46_in[415:384], zll_main_loop46_in[1765:1734], zll_main_loop46_in[517:486], zll_main_loop46_in[645:614], zll_main_loop46_in[479:448], zll_main_loop46_in[447:416], zll_main_loop46_in[1189:1158], zll_main_loop46_in[31:0], zll_main_loop46_in[2053:1798], zll_main_loop46_in[1157:646], zll_main_loop46_in[287:32], zll_main_loop46_in[485:480]};
  assign zll_main_loop96_in = {zll_main_loop116_in[2053:1542], zll_main_loop116_in[1541:1510], zll_main_loop116_in[1477:1446], zll_main_loop116_in[1445:1414], zll_main_loop116_in[1413:1382], zll_main_loop116_in[1381:1350], zll_main_loop116_in[1349:1318], zll_main_loop116_in[1317:1286], zll_main_loop116_in[1285:1254], zll_main_loop116_in[1253:1222], zll_main_loop116_in[1221:1190], zll_main_loop116_in[1189:1158], zll_main_loop116_in[1157:1126], zll_main_loop116_in[1125:1094], zll_main_loop116_in[1093:1062], zll_main_loop116_in[1061:1030], zll_main_loop116_in[1029:774], zll_main_loop116_in[773:262], zll_main_loop116_in[261:6], zll_main_loop116_in[5:0]};
  assign zll_main_loop_in = {zll_main_loop96_in[2021:1510], zll_main_loop96_in[1509:1478], zll_main_loop96_in[1445:1414], zll_main_loop96_in[1413:1382], zll_main_loop96_in[1381:1350], zll_main_loop96_in[1349:1318], zll_main_loop96_in[1317:1286], zll_main_loop96_in[1285:1254], zll_main_loop96_in[1253:1222], zll_main_loop96_in[1221:1190], zll_main_loop96_in[1189:1158], zll_main_loop96_in[1157:1126], zll_main_loop96_in[1125:1094], zll_main_loop96_in[1093:1062], zll_main_loop96_in[1061:1030], zll_main_loop96_in[1029:774], zll_main_loop96_in[773:262], zll_main_loop96_in[261:6], zll_main_loop96_in[5:0]};
  assign zll_main_loop38_in = {zll_main_loop_in[1989:1478], zll_main_loop_in[1477:1446], zll_main_loop_in[1413:1382], zll_main_loop_in[1381:1350], zll_main_loop_in[1349:1318], zll_main_loop_in[1317:1286], zll_main_loop_in[1285:1254], zll_main_loop_in[1253:1222], zll_main_loop_in[1221:1190], zll_main_loop_in[1189:1158], zll_main_loop_in[1157:1126], zll_main_loop_in[1125:1094], zll_main_loop_in[1093:1062], zll_main_loop_in[1061:1030], zll_main_loop_in[1029:774], zll_main_loop_in[773:262], zll_main_loop_in[261:6], zll_main_loop_in[5:0]};
  assign zll_main_loop54_in = {zll_main_loop38_in[1957:1446], zll_main_loop38_in[1445:1414], zll_main_loop38_in[1381:1350], zll_main_loop38_in[1349:1318], zll_main_loop38_in[1317:1286], zll_main_loop38_in[1285:1254], zll_main_loop38_in[1253:1222], zll_main_loop38_in[1221:1190], zll_main_loop38_in[1189:1158], zll_main_loop38_in[1157:1126], zll_main_loop38_in[1125:1094], zll_main_loop38_in[1093:1062], zll_main_loop38_in[1061:1030], zll_main_loop38_in[1029:774], zll_main_loop38_in[773:262], zll_main_loop38_in[261:6], zll_main_loop38_in[5:0]};
  assign zll_main_loop157_in = {zll_main_loop54_in[1925:1414], zll_main_loop54_in[1413:1382], zll_main_loop54_in[1349:1318], zll_main_loop54_in[1317:1286], zll_main_loop54_in[1285:1254], zll_main_loop54_in[1253:1222], zll_main_loop54_in[1221:1190], zll_main_loop54_in[1189:1158], zll_main_loop54_in[1157:1126], zll_main_loop54_in[1125:1094], zll_main_loop54_in[1093:1062], zll_main_loop54_in[1061:1030], zll_main_loop54_in[1029:774], zll_main_loop54_in[773:262], zll_main_loop54_in[261:6], zll_main_loop54_in[5:0]};
  assign zll_main_loop11_in = {zll_main_loop157_in[1893:1382], zll_main_loop157_in[1381:1350], zll_main_loop157_in[1317:1286], zll_main_loop157_in[1285:1254], zll_main_loop157_in[1253:1222], zll_main_loop157_in[1221:1190], zll_main_loop157_in[1189:1158], zll_main_loop157_in[1157:1126], zll_main_loop157_in[1125:1094], zll_main_loop157_in[1093:1062], zll_main_loop157_in[1061:1030], zll_main_loop157_in[1029:774], zll_main_loop157_in[773:262], zll_main_loop157_in[261:6], zll_main_loop157_in[5:0]};
  assign zll_main_loop132_in = {zll_main_loop11_in[1861:1350], zll_main_loop11_in[1349:1318], zll_main_loop11_in[1285:1254], zll_main_loop11_in[1253:1222], zll_main_loop11_in[1221:1190], zll_main_loop11_in[1189:1158], zll_main_loop11_in[1157:1126], zll_main_loop11_in[1125:1094], zll_main_loop11_in[1093:1062], zll_main_loop11_in[1061:1030], zll_main_loop11_in[1029:774], zll_main_loop11_in[773:262], zll_main_loop11_in[261:6], zll_main_loop11_in[5:0]};
  assign zll_main_loop77_in = {zll_main_loop132_in[1829:1318], zll_main_loop132_in[1317:1286], zll_main_loop132_in[1253:1222], zll_main_loop132_in[1221:1190], zll_main_loop132_in[1189:1158], zll_main_loop132_in[1157:1126], zll_main_loop132_in[1125:1094], zll_main_loop132_in[1093:1062], zll_main_loop132_in[1061:1030], zll_main_loop132_in[1029:774], zll_main_loop132_in[773:262], zll_main_loop132_in[261:6], zll_main_loop132_in[5:0]};
  assign zll_main_loop136_in = {zll_main_loop77_in[1797:1286], zll_main_loop77_in[1285:1254], zll_main_loop77_in[1221:1190], zll_main_loop77_in[1189:1158], zll_main_loop77_in[1157:1126], zll_main_loop77_in[1125:1094], zll_main_loop77_in[1093:1062], zll_main_loop77_in[1061:1030], zll_main_loop77_in[1029:774], zll_main_loop77_in[773:262], zll_main_loop77_in[261:6], zll_main_loop77_in[5:0]};
  assign zll_main_loop150_in = {zll_main_loop136_in[1765:1254], zll_main_loop136_in[1253:1222], zll_main_loop136_in[1189:1158], zll_main_loop136_in[1157:1126], zll_main_loop136_in[1125:1094], zll_main_loop136_in[1093:1062], zll_main_loop136_in[1061:1030], zll_main_loop136_in[1029:774], zll_main_loop136_in[773:262], zll_main_loop136_in[261:6], zll_main_loop136_in[5:0]};
  assign zll_main_loop75_in = {zll_main_loop150_in[1733:1222], zll_main_loop150_in[1221:1190], zll_main_loop150_in[1157:1126], zll_main_loop150_in[1125:1094], zll_main_loop150_in[1093:1062], zll_main_loop150_in[1061:1030], zll_main_loop150_in[1029:774], zll_main_loop150_in[773:262], zll_main_loop150_in[261:6], zll_main_loop150_in[5:0]};
  assign zll_main_loop19_in = {zll_main_loop75_in[1701:1190], zll_main_loop75_in[1189:1158], zll_main_loop75_in[1125:1094], zll_main_loop75_in[1093:1062], zll_main_loop75_in[1061:1030], zll_main_loop75_in[1029:774], zll_main_loop75_in[773:262], zll_main_loop75_in[261:6], zll_main_loop75_in[5:0]};
  assign zll_main_loop146_in = {zll_main_loop19_in[1669:1158], zll_main_loop19_in[1157:1126], zll_main_loop19_in[1093:1062], zll_main_loop19_in[1061:1030], zll_main_loop19_in[1029:774], zll_main_loop19_in[773:262], zll_main_loop19_in[261:6], zll_main_loop19_in[5:0]};
  assign zll_main_loop141_in = {zll_main_loop146_in[1637:1126], zll_main_loop146_in[1125:1094], zll_main_loop146_in[1061:1030], zll_main_loop146_in[1029:774], zll_main_loop146_in[773:262], zll_main_loop146_in[261:6], zll_main_loop146_in[5:0]};
  assign main_updatesched_in = zll_main_loop141_in[1605:1094];
  assign zll_main_updatesched4_in = main_updatesched_in[511:0];
  assign zll_main_updatesched13_in = {zll_main_updatesched4_in[479:448], zll_main_updatesched4_in[511:480], zll_main_updatesched4_in[447:416], zll_main_updatesched4_in[415:384], zll_main_updatesched4_in[383:352], zll_main_updatesched4_in[351:320], zll_main_updatesched4_in[319:288], zll_main_updatesched4_in[287:256], zll_main_updatesched4_in[255:224], zll_main_updatesched4_in[223:192], zll_main_updatesched4_in[191:160], zll_main_updatesched4_in[159:128], zll_main_updatesched4_in[127:96], zll_main_updatesched4_in[95:64], zll_main_updatesched4_in[63:32], zll_main_updatesched4_in[31:0]};
  assign zll_main_updatesched3_in = {zll_main_updatesched13_in[447:416], zll_main_updatesched13_in[511:480], zll_main_updatesched13_in[479:448], zll_main_updatesched13_in[415:384], zll_main_updatesched13_in[383:352], zll_main_updatesched13_in[351:320], zll_main_updatesched13_in[319:288], zll_main_updatesched13_in[287:256], zll_main_updatesched13_in[255:224], zll_main_updatesched13_in[223:192], zll_main_updatesched13_in[191:160], zll_main_updatesched13_in[159:128], zll_main_updatesched13_in[127:96], zll_main_updatesched13_in[95:64], zll_main_updatesched13_in[63:32], zll_main_updatesched13_in[31:0]};
  assign zll_main_updatesched15_in = {zll_main_updatesched3_in[511:480], zll_main_updatesched3_in[479:448], zll_main_updatesched3_in[415:384], zll_main_updatesched3_in[447:416], zll_main_updatesched3_in[383:352], zll_main_updatesched3_in[351:320], zll_main_updatesched3_in[319:288], zll_main_updatesched3_in[287:256], zll_main_updatesched3_in[255:224], zll_main_updatesched3_in[223:192], zll_main_updatesched3_in[191:160], zll_main_updatesched3_in[159:128], zll_main_updatesched3_in[127:96], zll_main_updatesched3_in[95:64], zll_main_updatesched3_in[63:32], zll_main_updatesched3_in[31:0]};
  assign zll_main_updatesched7_in = {zll_main_updatesched15_in[511:480], zll_main_updatesched15_in[479:448], zll_main_updatesched15_in[447:416], zll_main_updatesched15_in[351:320], zll_main_updatesched15_in[415:384], zll_main_updatesched15_in[383:352], zll_main_updatesched15_in[319:288], zll_main_updatesched15_in[287:256], zll_main_updatesched15_in[255:224], zll_main_updatesched15_in[223:192], zll_main_updatesched15_in[191:160], zll_main_updatesched15_in[159:128], zll_main_updatesched15_in[127:96], zll_main_updatesched15_in[95:64], zll_main_updatesched15_in[63:32], zll_main_updatesched15_in[31:0]};
  assign zll_main_updatesched5_in = {zll_main_updatesched7_in[511:480], zll_main_updatesched7_in[479:448], zll_main_updatesched7_in[447:416], zll_main_updatesched7_in[415:384], zll_main_updatesched7_in[319:288], zll_main_updatesched7_in[383:352], zll_main_updatesched7_in[351:320], zll_main_updatesched7_in[287:256], zll_main_updatesched7_in[255:224], zll_main_updatesched7_in[223:192], zll_main_updatesched7_in[191:160], zll_main_updatesched7_in[159:128], zll_main_updatesched7_in[127:96], zll_main_updatesched7_in[95:64], zll_main_updatesched7_in[63:32], zll_main_updatesched7_in[31:0]};
  assign zll_main_updatesched_in = {zll_main_updatesched5_in[287:256], zll_main_updatesched5_in[511:480], zll_main_updatesched5_in[479:448], zll_main_updatesched5_in[447:416], zll_main_updatesched5_in[415:384], zll_main_updatesched5_in[383:352], zll_main_updatesched5_in[351:320], zll_main_updatesched5_in[319:288], zll_main_updatesched5_in[255:224], zll_main_updatesched5_in[223:192], zll_main_updatesched5_in[191:160], zll_main_updatesched5_in[159:128], zll_main_updatesched5_in[127:96], zll_main_updatesched5_in[95:64], zll_main_updatesched5_in[63:32], zll_main_updatesched5_in[31:0]};
  assign zll_main_updatesched1_in = {zll_main_updatesched_in[511:480], zll_main_updatesched_in[479:448], zll_main_updatesched_in[447:416], zll_main_updatesched_in[415:384], zll_main_updatesched_in[383:352], zll_main_updatesched_in[351:320], zll_main_updatesched_in[319:288], zll_main_updatesched_in[255:224], zll_main_updatesched_in[287:256], zll_main_updatesched_in[223:192], zll_main_updatesched_in[191:160], zll_main_updatesched_in[159:128], zll_main_updatesched_in[127:96], zll_main_updatesched_in[95:64], zll_main_updatesched_in[63:32], zll_main_updatesched_in[31:0]};
  assign zll_main_updatesched6_in = {zll_main_updatesched1_in[511:480], zll_main_updatesched1_in[479:448], zll_main_updatesched1_in[223:192], zll_main_updatesched1_in[447:416], zll_main_updatesched1_in[415:384], zll_main_updatesched1_in[383:352], zll_main_updatesched1_in[351:320], zll_main_updatesched1_in[319:288], zll_main_updatesched1_in[287:256], zll_main_updatesched1_in[255:224], zll_main_updatesched1_in[191:160], zll_main_updatesched1_in[159:128], zll_main_updatesched1_in[127:96], zll_main_updatesched1_in[95:64], zll_main_updatesched1_in[63:32], zll_main_updatesched1_in[31:0]};
  assign zll_main_updatesched8_in = {zll_main_updatesched6_in[191:160], zll_main_updatesched6_in[511:480], zll_main_updatesched6_in[479:448], zll_main_updatesched6_in[447:416], zll_main_updatesched6_in[415:384], zll_main_updatesched6_in[383:352], zll_main_updatesched6_in[351:320], zll_main_updatesched6_in[319:288], zll_main_updatesched6_in[287:256], zll_main_updatesched6_in[255:224], zll_main_updatesched6_in[223:192], zll_main_updatesched6_in[159:128], zll_main_updatesched6_in[127:96], zll_main_updatesched6_in[95:64], zll_main_updatesched6_in[63:32], zll_main_updatesched6_in[31:0]};
  assign zll_main_updatesched12_in = {zll_main_updatesched8_in[511:480], zll_main_updatesched8_in[479:448], zll_main_updatesched8_in[447:416], zll_main_updatesched8_in[415:384], zll_main_updatesched8_in[383:352], zll_main_updatesched8_in[351:320], zll_main_updatesched8_in[319:288], zll_main_updatesched8_in[159:128], zll_main_updatesched8_in[287:256], zll_main_updatesched8_in[255:224], zll_main_updatesched8_in[223:192], zll_main_updatesched8_in[191:160], zll_main_updatesched8_in[127:96], zll_main_updatesched8_in[95:64], zll_main_updatesched8_in[63:32], zll_main_updatesched8_in[31:0]};
  assign zll_main_updatesched14_in = {zll_main_updatesched12_in[511:480], zll_main_updatesched12_in[479:448], zll_main_updatesched12_in[447:416], zll_main_updatesched12_in[415:384], zll_main_updatesched12_in[383:352], zll_main_updatesched12_in[351:320], zll_main_updatesched12_in[319:288], zll_main_updatesched12_in[127:96], zll_main_updatesched12_in[287:256], zll_main_updatesched12_in[255:224], zll_main_updatesched12_in[223:192], zll_main_updatesched12_in[191:160], zll_main_updatesched12_in[159:128], zll_main_updatesched12_in[95:64], zll_main_updatesched12_in[63:32], zll_main_updatesched12_in[31:0]};
  assign zll_main_updatesched2_in = {zll_main_updatesched14_in[511:480], zll_main_updatesched14_in[479:448], zll_main_updatesched14_in[447:416], zll_main_updatesched14_in[415:384], zll_main_updatesched14_in[383:352], zll_main_updatesched14_in[95:64], zll_main_updatesched14_in[351:320], zll_main_updatesched14_in[319:288], zll_main_updatesched14_in[287:256], zll_main_updatesched14_in[255:224], zll_main_updatesched14_in[223:192], zll_main_updatesched14_in[191:160], zll_main_updatesched14_in[159:128], zll_main_updatesched14_in[127:96], zll_main_updatesched14_in[63:32], zll_main_updatesched14_in[31:0]};
  assign main_sigma1_in = zll_main_updatesched2_in[63:32];
  assign main_rotater17_in = main_sigma1_in[31:0];
  assign zll_main_rotater1729_in = main_rotater17_in[31:0];
  assign zll_main_rotater1710_in = {zll_main_rotater1729_in[31], zll_main_rotater1729_in[29], zll_main_rotater1729_in[30], zll_main_rotater1729_in[28], zll_main_rotater1729_in[27], zll_main_rotater1729_in[26], zll_main_rotater1729_in[25], zll_main_rotater1729_in[24], zll_main_rotater1729_in[23], zll_main_rotater1729_in[22], zll_main_rotater1729_in[21], zll_main_rotater1729_in[20], zll_main_rotater1729_in[19], zll_main_rotater1729_in[18], zll_main_rotater1729_in[17], zll_main_rotater1729_in[16], zll_main_rotater1729_in[15], zll_main_rotater1729_in[14], zll_main_rotater1729_in[13], zll_main_rotater1729_in[12], zll_main_rotater1729_in[11], zll_main_rotater1729_in[10], zll_main_rotater1729_in[9], zll_main_rotater1729_in[8], zll_main_rotater1729_in[7], zll_main_rotater1729_in[6], zll_main_rotater1729_in[5], zll_main_rotater1729_in[4], zll_main_rotater1729_in[3], zll_main_rotater1729_in[2], zll_main_rotater1729_in[1], zll_main_rotater1729_in[0]};
  assign zll_main_rotater1727_in = {zll_main_rotater1710_in[31], zll_main_rotater1710_in[28], zll_main_rotater1710_in[30], zll_main_rotater1710_in[29], zll_main_rotater1710_in[27], zll_main_rotater1710_in[26], zll_main_rotater1710_in[25], zll_main_rotater1710_in[24], zll_main_rotater1710_in[23], zll_main_rotater1710_in[22], zll_main_rotater1710_in[21], zll_main_rotater1710_in[20], zll_main_rotater1710_in[19], zll_main_rotater1710_in[18], zll_main_rotater1710_in[17], zll_main_rotater1710_in[16], zll_main_rotater1710_in[15], zll_main_rotater1710_in[14], zll_main_rotater1710_in[13], zll_main_rotater1710_in[12], zll_main_rotater1710_in[11], zll_main_rotater1710_in[10], zll_main_rotater1710_in[9], zll_main_rotater1710_in[8], zll_main_rotater1710_in[7], zll_main_rotater1710_in[6], zll_main_rotater1710_in[5], zll_main_rotater1710_in[4], zll_main_rotater1710_in[3], zll_main_rotater1710_in[2], zll_main_rotater1710_in[1], zll_main_rotater1710_in[0]};
  assign zll_main_rotater1724_in = {zll_main_rotater1727_in[31], zll_main_rotater1727_in[30], zll_main_rotater1727_in[27], zll_main_rotater1727_in[29], zll_main_rotater1727_in[28], zll_main_rotater1727_in[26], zll_main_rotater1727_in[25], zll_main_rotater1727_in[24], zll_main_rotater1727_in[23], zll_main_rotater1727_in[22], zll_main_rotater1727_in[21], zll_main_rotater1727_in[20], zll_main_rotater1727_in[19], zll_main_rotater1727_in[18], zll_main_rotater1727_in[17], zll_main_rotater1727_in[16], zll_main_rotater1727_in[15], zll_main_rotater1727_in[14], zll_main_rotater1727_in[13], zll_main_rotater1727_in[12], zll_main_rotater1727_in[11], zll_main_rotater1727_in[10], zll_main_rotater1727_in[9], zll_main_rotater1727_in[8], zll_main_rotater1727_in[7], zll_main_rotater1727_in[6], zll_main_rotater1727_in[5], zll_main_rotater1727_in[4], zll_main_rotater1727_in[3], zll_main_rotater1727_in[2], zll_main_rotater1727_in[1], zll_main_rotater1727_in[0]};
  assign zll_main_rotater1730_in = {zll_main_rotater1724_in[31], zll_main_rotater1724_in[30], zll_main_rotater1724_in[29], zll_main_rotater1724_in[26], zll_main_rotater1724_in[28], zll_main_rotater1724_in[27], zll_main_rotater1724_in[25], zll_main_rotater1724_in[24], zll_main_rotater1724_in[23], zll_main_rotater1724_in[22], zll_main_rotater1724_in[21], zll_main_rotater1724_in[20], zll_main_rotater1724_in[19], zll_main_rotater1724_in[18], zll_main_rotater1724_in[17], zll_main_rotater1724_in[16], zll_main_rotater1724_in[15], zll_main_rotater1724_in[14], zll_main_rotater1724_in[13], zll_main_rotater1724_in[12], zll_main_rotater1724_in[11], zll_main_rotater1724_in[10], zll_main_rotater1724_in[9], zll_main_rotater1724_in[8], zll_main_rotater1724_in[7], zll_main_rotater1724_in[6], zll_main_rotater1724_in[5], zll_main_rotater1724_in[4], zll_main_rotater1724_in[3], zll_main_rotater1724_in[2], zll_main_rotater1724_in[1], zll_main_rotater1724_in[0]};
  assign zll_main_rotater178_in = {zll_main_rotater1730_in[31], zll_main_rotater1730_in[30], zll_main_rotater1730_in[29], zll_main_rotater1730_in[28], zll_main_rotater1730_in[27], zll_main_rotater1730_in[26], zll_main_rotater1730_in[24], zll_main_rotater1730_in[25], zll_main_rotater1730_in[23], zll_main_rotater1730_in[22], zll_main_rotater1730_in[21], zll_main_rotater1730_in[20], zll_main_rotater1730_in[19], zll_main_rotater1730_in[18], zll_main_rotater1730_in[17], zll_main_rotater1730_in[16], zll_main_rotater1730_in[15], zll_main_rotater1730_in[14], zll_main_rotater1730_in[13], zll_main_rotater1730_in[12], zll_main_rotater1730_in[11], zll_main_rotater1730_in[10], zll_main_rotater1730_in[9], zll_main_rotater1730_in[8], zll_main_rotater1730_in[7], zll_main_rotater1730_in[6], zll_main_rotater1730_in[5], zll_main_rotater1730_in[4], zll_main_rotater1730_in[3], zll_main_rotater1730_in[2], zll_main_rotater1730_in[1], zll_main_rotater1730_in[0]};
  assign zll_main_rotater177_in = {zll_main_rotater178_in[31], zll_main_rotater178_in[30], zll_main_rotater178_in[29], zll_main_rotater178_in[22], zll_main_rotater178_in[28], zll_main_rotater178_in[27], zll_main_rotater178_in[26], zll_main_rotater178_in[25], zll_main_rotater178_in[24], zll_main_rotater178_in[23], zll_main_rotater178_in[21], zll_main_rotater178_in[20], zll_main_rotater178_in[19], zll_main_rotater178_in[18], zll_main_rotater178_in[17], zll_main_rotater178_in[16], zll_main_rotater178_in[15], zll_main_rotater178_in[14], zll_main_rotater178_in[13], zll_main_rotater178_in[12], zll_main_rotater178_in[11], zll_main_rotater178_in[10], zll_main_rotater178_in[9], zll_main_rotater178_in[8], zll_main_rotater178_in[7], zll_main_rotater178_in[6], zll_main_rotater178_in[5], zll_main_rotater178_in[4], zll_main_rotater178_in[3], zll_main_rotater178_in[2], zll_main_rotater178_in[1], zll_main_rotater178_in[0]};
  assign zll_main_rotater175_in = {zll_main_rotater177_in[31], zll_main_rotater177_in[30], zll_main_rotater177_in[29], zll_main_rotater177_in[28], zll_main_rotater177_in[27], zll_main_rotater177_in[26], zll_main_rotater177_in[21], zll_main_rotater177_in[25], zll_main_rotater177_in[24], zll_main_rotater177_in[23], zll_main_rotater177_in[22], zll_main_rotater177_in[20], zll_main_rotater177_in[19], zll_main_rotater177_in[18], zll_main_rotater177_in[17], zll_main_rotater177_in[16], zll_main_rotater177_in[15], zll_main_rotater177_in[14], zll_main_rotater177_in[13], zll_main_rotater177_in[12], zll_main_rotater177_in[11], zll_main_rotater177_in[10], zll_main_rotater177_in[9], zll_main_rotater177_in[8], zll_main_rotater177_in[7], zll_main_rotater177_in[6], zll_main_rotater177_in[5], zll_main_rotater177_in[4], zll_main_rotater177_in[3], zll_main_rotater177_in[2], zll_main_rotater177_in[1], zll_main_rotater177_in[0]};
  assign zll_main_rotater1714_in = {zll_main_rotater175_in[31], zll_main_rotater175_in[30], zll_main_rotater175_in[20], zll_main_rotater175_in[29], zll_main_rotater175_in[28], zll_main_rotater175_in[27], zll_main_rotater175_in[26], zll_main_rotater175_in[25], zll_main_rotater175_in[24], zll_main_rotater175_in[23], zll_main_rotater175_in[22], zll_main_rotater175_in[21], zll_main_rotater175_in[19], zll_main_rotater175_in[18], zll_main_rotater175_in[17], zll_main_rotater175_in[16], zll_main_rotater175_in[15], zll_main_rotater175_in[14], zll_main_rotater175_in[13], zll_main_rotater175_in[12], zll_main_rotater175_in[11], zll_main_rotater175_in[10], zll_main_rotater175_in[9], zll_main_rotater175_in[8], zll_main_rotater175_in[7], zll_main_rotater175_in[6], zll_main_rotater175_in[5], zll_main_rotater175_in[4], zll_main_rotater175_in[3], zll_main_rotater175_in[2], zll_main_rotater175_in[1], zll_main_rotater175_in[0]};
  assign zll_main_rotater1721_in = {zll_main_rotater1714_in[31], zll_main_rotater1714_in[30], zll_main_rotater1714_in[29], zll_main_rotater1714_in[28], zll_main_rotater1714_in[18], zll_main_rotater1714_in[27], zll_main_rotater1714_in[26], zll_main_rotater1714_in[25], zll_main_rotater1714_in[24], zll_main_rotater1714_in[23], zll_main_rotater1714_in[22], zll_main_rotater1714_in[21], zll_main_rotater1714_in[20], zll_main_rotater1714_in[19], zll_main_rotater1714_in[17], zll_main_rotater1714_in[16], zll_main_rotater1714_in[15], zll_main_rotater1714_in[14], zll_main_rotater1714_in[13], zll_main_rotater1714_in[12], zll_main_rotater1714_in[11], zll_main_rotater1714_in[10], zll_main_rotater1714_in[9], zll_main_rotater1714_in[8], zll_main_rotater1714_in[7], zll_main_rotater1714_in[6], zll_main_rotater1714_in[5], zll_main_rotater1714_in[4], zll_main_rotater1714_in[3], zll_main_rotater1714_in[2], zll_main_rotater1714_in[1], zll_main_rotater1714_in[0]};
  assign zll_main_rotater1712_in = {zll_main_rotater1721_in[31], zll_main_rotater1721_in[30], zll_main_rotater1721_in[29], zll_main_rotater1721_in[28], zll_main_rotater1721_in[27], zll_main_rotater1721_in[26], zll_main_rotater1721_in[25], zll_main_rotater1721_in[24], zll_main_rotater1721_in[23], zll_main_rotater1721_in[22], zll_main_rotater1721_in[17], zll_main_rotater1721_in[21], zll_main_rotater1721_in[20], zll_main_rotater1721_in[19], zll_main_rotater1721_in[18], zll_main_rotater1721_in[16], zll_main_rotater1721_in[15], zll_main_rotater1721_in[14], zll_main_rotater1721_in[13], zll_main_rotater1721_in[12], zll_main_rotater1721_in[11], zll_main_rotater1721_in[10], zll_main_rotater1721_in[9], zll_main_rotater1721_in[8], zll_main_rotater1721_in[7], zll_main_rotater1721_in[6], zll_main_rotater1721_in[5], zll_main_rotater1721_in[4], zll_main_rotater1721_in[3], zll_main_rotater1721_in[2], zll_main_rotater1721_in[1], zll_main_rotater1721_in[0]};
  assign zll_main_rotater171_in = {zll_main_rotater1712_in[31], zll_main_rotater1712_in[30], zll_main_rotater1712_in[29], zll_main_rotater1712_in[28], zll_main_rotater1712_in[27], zll_main_rotater1712_in[26], zll_main_rotater1712_in[25], zll_main_rotater1712_in[24], zll_main_rotater1712_in[23], zll_main_rotater1712_in[22], zll_main_rotater1712_in[21], zll_main_rotater1712_in[20], zll_main_rotater1712_in[16], zll_main_rotater1712_in[19], zll_main_rotater1712_in[18], zll_main_rotater1712_in[17], zll_main_rotater1712_in[15], zll_main_rotater1712_in[14], zll_main_rotater1712_in[13], zll_main_rotater1712_in[12], zll_main_rotater1712_in[11], zll_main_rotater1712_in[10], zll_main_rotater1712_in[9], zll_main_rotater1712_in[8], zll_main_rotater1712_in[7], zll_main_rotater1712_in[6], zll_main_rotater1712_in[5], zll_main_rotater1712_in[4], zll_main_rotater1712_in[3], zll_main_rotater1712_in[2], zll_main_rotater1712_in[1], zll_main_rotater1712_in[0]};
  assign zll_main_rotater1711_in = {zll_main_rotater171_in[31], zll_main_rotater171_in[30], zll_main_rotater171_in[29], zll_main_rotater171_in[28], zll_main_rotater171_in[27], zll_main_rotater171_in[26], zll_main_rotater171_in[25], zll_main_rotater171_in[24], zll_main_rotater171_in[23], zll_main_rotater171_in[22], zll_main_rotater171_in[15], zll_main_rotater171_in[21], zll_main_rotater171_in[20], zll_main_rotater171_in[19], zll_main_rotater171_in[18], zll_main_rotater171_in[17], zll_main_rotater171_in[16], zll_main_rotater171_in[14], zll_main_rotater171_in[13], zll_main_rotater171_in[12], zll_main_rotater171_in[11], zll_main_rotater171_in[10], zll_main_rotater171_in[9], zll_main_rotater171_in[8], zll_main_rotater171_in[7], zll_main_rotater171_in[6], zll_main_rotater171_in[5], zll_main_rotater171_in[4], zll_main_rotater171_in[3], zll_main_rotater171_in[2], zll_main_rotater171_in[1], zll_main_rotater171_in[0]};
  assign zll_main_rotater1723_in = {zll_main_rotater1711_in[31], zll_main_rotater1711_in[30], zll_main_rotater1711_in[29], zll_main_rotater1711_in[14], zll_main_rotater1711_in[28], zll_main_rotater1711_in[27], zll_main_rotater1711_in[26], zll_main_rotater1711_in[25], zll_main_rotater1711_in[24], zll_main_rotater1711_in[23], zll_main_rotater1711_in[22], zll_main_rotater1711_in[21], zll_main_rotater1711_in[20], zll_main_rotater1711_in[19], zll_main_rotater1711_in[18], zll_main_rotater1711_in[17], zll_main_rotater1711_in[16], zll_main_rotater1711_in[15], zll_main_rotater1711_in[13], zll_main_rotater1711_in[12], zll_main_rotater1711_in[11], zll_main_rotater1711_in[10], zll_main_rotater1711_in[9], zll_main_rotater1711_in[8], zll_main_rotater1711_in[7], zll_main_rotater1711_in[6], zll_main_rotater1711_in[5], zll_main_rotater1711_in[4], zll_main_rotater1711_in[3], zll_main_rotater1711_in[2], zll_main_rotater1711_in[1], zll_main_rotater1711_in[0]};
  assign zll_main_rotater1717_in = {zll_main_rotater1723_in[31], zll_main_rotater1723_in[30], zll_main_rotater1723_in[29], zll_main_rotater1723_in[28], zll_main_rotater1723_in[27], zll_main_rotater1723_in[26], zll_main_rotater1723_in[25], zll_main_rotater1723_in[24], zll_main_rotater1723_in[23], zll_main_rotater1723_in[22], zll_main_rotater1723_in[21], zll_main_rotater1723_in[20], zll_main_rotater1723_in[19], zll_main_rotater1723_in[18], zll_main_rotater1723_in[17], zll_main_rotater1723_in[16], zll_main_rotater1723_in[13], zll_main_rotater1723_in[15], zll_main_rotater1723_in[14], zll_main_rotater1723_in[12], zll_main_rotater1723_in[11], zll_main_rotater1723_in[10], zll_main_rotater1723_in[9], zll_main_rotater1723_in[8], zll_main_rotater1723_in[7], zll_main_rotater1723_in[6], zll_main_rotater1723_in[5], zll_main_rotater1723_in[4], zll_main_rotater1723_in[3], zll_main_rotater1723_in[2], zll_main_rotater1723_in[1], zll_main_rotater1723_in[0]};
  assign zll_main_rotater1715_in = {zll_main_rotater1717_in[31], zll_main_rotater1717_in[30], zll_main_rotater1717_in[29], zll_main_rotater1717_in[28], zll_main_rotater1717_in[27], zll_main_rotater1717_in[26], zll_main_rotater1717_in[25], zll_main_rotater1717_in[24], zll_main_rotater1717_in[23], zll_main_rotater1717_in[22], zll_main_rotater1717_in[21], zll_main_rotater1717_in[20], zll_main_rotater1717_in[11], zll_main_rotater1717_in[19], zll_main_rotater1717_in[18], zll_main_rotater1717_in[17], zll_main_rotater1717_in[16], zll_main_rotater1717_in[15], zll_main_rotater1717_in[14], zll_main_rotater1717_in[13], zll_main_rotater1717_in[12], zll_main_rotater1717_in[10], zll_main_rotater1717_in[9], zll_main_rotater1717_in[8], zll_main_rotater1717_in[7], zll_main_rotater1717_in[6], zll_main_rotater1717_in[5], zll_main_rotater1717_in[4], zll_main_rotater1717_in[3], zll_main_rotater1717_in[2], zll_main_rotater1717_in[1], zll_main_rotater1717_in[0]};
  assign zll_main_rotater1716_in = {zll_main_rotater1715_in[31], zll_main_rotater1715_in[30], zll_main_rotater1715_in[29], zll_main_rotater1715_in[28], zll_main_rotater1715_in[27], zll_main_rotater1715_in[26], zll_main_rotater1715_in[25], zll_main_rotater1715_in[24], zll_main_rotater1715_in[23], zll_main_rotater1715_in[22], zll_main_rotater1715_in[21], zll_main_rotater1715_in[20], zll_main_rotater1715_in[19], zll_main_rotater1715_in[18], zll_main_rotater1715_in[17], zll_main_rotater1715_in[10], zll_main_rotater1715_in[16], zll_main_rotater1715_in[15], zll_main_rotater1715_in[14], zll_main_rotater1715_in[13], zll_main_rotater1715_in[12], zll_main_rotater1715_in[11], zll_main_rotater1715_in[9], zll_main_rotater1715_in[8], zll_main_rotater1715_in[7], zll_main_rotater1715_in[6], zll_main_rotater1715_in[5], zll_main_rotater1715_in[4], zll_main_rotater1715_in[3], zll_main_rotater1715_in[2], zll_main_rotater1715_in[1], zll_main_rotater1715_in[0]};
  assign zll_main_rotater179_in = {zll_main_rotater1716_in[31], zll_main_rotater1716_in[30], zll_main_rotater1716_in[29], zll_main_rotater1716_in[28], zll_main_rotater1716_in[27], zll_main_rotater1716_in[26], zll_main_rotater1716_in[25], zll_main_rotater1716_in[24], zll_main_rotater1716_in[23], zll_main_rotater1716_in[22], zll_main_rotater1716_in[21], zll_main_rotater1716_in[20], zll_main_rotater1716_in[19], zll_main_rotater1716_in[18], zll_main_rotater1716_in[17], zll_main_rotater1716_in[9], zll_main_rotater1716_in[16], zll_main_rotater1716_in[15], zll_main_rotater1716_in[14], zll_main_rotater1716_in[13], zll_main_rotater1716_in[12], zll_main_rotater1716_in[11], zll_main_rotater1716_in[10], zll_main_rotater1716_in[8], zll_main_rotater1716_in[7], zll_main_rotater1716_in[6], zll_main_rotater1716_in[5], zll_main_rotater1716_in[4], zll_main_rotater1716_in[3], zll_main_rotater1716_in[2], zll_main_rotater1716_in[1], zll_main_rotater1716_in[0]};
  assign zll_main_rotater173_in = {zll_main_rotater179_in[31], zll_main_rotater179_in[30], zll_main_rotater179_in[29], zll_main_rotater179_in[28], zll_main_rotater179_in[8], zll_main_rotater179_in[27], zll_main_rotater179_in[26], zll_main_rotater179_in[25], zll_main_rotater179_in[24], zll_main_rotater179_in[23], zll_main_rotater179_in[22], zll_main_rotater179_in[21], zll_main_rotater179_in[20], zll_main_rotater179_in[19], zll_main_rotater179_in[18], zll_main_rotater179_in[17], zll_main_rotater179_in[16], zll_main_rotater179_in[15], zll_main_rotater179_in[14], zll_main_rotater179_in[13], zll_main_rotater179_in[12], zll_main_rotater179_in[11], zll_main_rotater179_in[10], zll_main_rotater179_in[9], zll_main_rotater179_in[7], zll_main_rotater179_in[6], zll_main_rotater179_in[5], zll_main_rotater179_in[4], zll_main_rotater179_in[3], zll_main_rotater179_in[2], zll_main_rotater179_in[1], zll_main_rotater179_in[0]};
  assign zll_main_rotater1726_in = {zll_main_rotater173_in[31], zll_main_rotater173_in[30], zll_main_rotater173_in[29], zll_main_rotater173_in[28], zll_main_rotater173_in[27], zll_main_rotater173_in[26], zll_main_rotater173_in[25], zll_main_rotater173_in[24], zll_main_rotater173_in[23], zll_main_rotater173_in[22], zll_main_rotater173_in[21], zll_main_rotater173_in[20], zll_main_rotater173_in[19], zll_main_rotater173_in[18], zll_main_rotater173_in[17], zll_main_rotater173_in[16], zll_main_rotater173_in[15], zll_main_rotater173_in[14], zll_main_rotater173_in[13], zll_main_rotater173_in[7], zll_main_rotater173_in[12], zll_main_rotater173_in[11], zll_main_rotater173_in[10], zll_main_rotater173_in[9], zll_main_rotater173_in[8], zll_main_rotater173_in[6], zll_main_rotater173_in[5], zll_main_rotater173_in[4], zll_main_rotater173_in[3], zll_main_rotater173_in[2], zll_main_rotater173_in[1], zll_main_rotater173_in[0]};
  assign zll_main_rotater176_in = {zll_main_rotater1726_in[31], zll_main_rotater1726_in[30], zll_main_rotater1726_in[29], zll_main_rotater1726_in[28], zll_main_rotater1726_in[27], zll_main_rotater1726_in[26], zll_main_rotater1726_in[25], zll_main_rotater1726_in[24], zll_main_rotater1726_in[23], zll_main_rotater1726_in[22], zll_main_rotater1726_in[21], zll_main_rotater1726_in[6], zll_main_rotater1726_in[20], zll_main_rotater1726_in[19], zll_main_rotater1726_in[18], zll_main_rotater1726_in[17], zll_main_rotater1726_in[16], zll_main_rotater1726_in[15], zll_main_rotater1726_in[14], zll_main_rotater1726_in[13], zll_main_rotater1726_in[12], zll_main_rotater1726_in[11], zll_main_rotater1726_in[10], zll_main_rotater1726_in[9], zll_main_rotater1726_in[8], zll_main_rotater1726_in[7], zll_main_rotater1726_in[5], zll_main_rotater1726_in[4], zll_main_rotater1726_in[3], zll_main_rotater1726_in[2], zll_main_rotater1726_in[1], zll_main_rotater1726_in[0]};
  assign zll_main_rotater1713_in = {zll_main_rotater176_in[31], zll_main_rotater176_in[30], zll_main_rotater176_in[29], zll_main_rotater176_in[28], zll_main_rotater176_in[27], zll_main_rotater176_in[26], zll_main_rotater176_in[25], zll_main_rotater176_in[24], zll_main_rotater176_in[23], zll_main_rotater176_in[22], zll_main_rotater176_in[21], zll_main_rotater176_in[20], zll_main_rotater176_in[19], zll_main_rotater176_in[18], zll_main_rotater176_in[17], zll_main_rotater176_in[5], zll_main_rotater176_in[16], zll_main_rotater176_in[15], zll_main_rotater176_in[14], zll_main_rotater176_in[13], zll_main_rotater176_in[12], zll_main_rotater176_in[11], zll_main_rotater176_in[10], zll_main_rotater176_in[9], zll_main_rotater176_in[8], zll_main_rotater176_in[7], zll_main_rotater176_in[6], zll_main_rotater176_in[4], zll_main_rotater176_in[3], zll_main_rotater176_in[2], zll_main_rotater176_in[1], zll_main_rotater176_in[0]};
  assign zll_main_rotater1728_in = {zll_main_rotater1713_in[31], zll_main_rotater1713_in[30], zll_main_rotater1713_in[29], zll_main_rotater1713_in[28], zll_main_rotater1713_in[27], zll_main_rotater1713_in[26], zll_main_rotater1713_in[25], zll_main_rotater1713_in[4], zll_main_rotater1713_in[24], zll_main_rotater1713_in[23], zll_main_rotater1713_in[22], zll_main_rotater1713_in[21], zll_main_rotater1713_in[20], zll_main_rotater1713_in[19], zll_main_rotater1713_in[18], zll_main_rotater1713_in[17], zll_main_rotater1713_in[16], zll_main_rotater1713_in[15], zll_main_rotater1713_in[14], zll_main_rotater1713_in[13], zll_main_rotater1713_in[12], zll_main_rotater1713_in[11], zll_main_rotater1713_in[10], zll_main_rotater1713_in[9], zll_main_rotater1713_in[8], zll_main_rotater1713_in[7], zll_main_rotater1713_in[6], zll_main_rotater1713_in[5], zll_main_rotater1713_in[3], zll_main_rotater1713_in[2], zll_main_rotater1713_in[1], zll_main_rotater1713_in[0]};
  assign zll_main_rotater17_in = {zll_main_rotater1728_in[31], zll_main_rotater1728_in[3], zll_main_rotater1728_in[30], zll_main_rotater1728_in[29], zll_main_rotater1728_in[28], zll_main_rotater1728_in[27], zll_main_rotater1728_in[26], zll_main_rotater1728_in[25], zll_main_rotater1728_in[24], zll_main_rotater1728_in[23], zll_main_rotater1728_in[22], zll_main_rotater1728_in[21], zll_main_rotater1728_in[20], zll_main_rotater1728_in[19], zll_main_rotater1728_in[18], zll_main_rotater1728_in[17], zll_main_rotater1728_in[16], zll_main_rotater1728_in[15], zll_main_rotater1728_in[14], zll_main_rotater1728_in[13], zll_main_rotater1728_in[12], zll_main_rotater1728_in[11], zll_main_rotater1728_in[10], zll_main_rotater1728_in[9], zll_main_rotater1728_in[8], zll_main_rotater1728_in[7], zll_main_rotater1728_in[6], zll_main_rotater1728_in[5], zll_main_rotater1728_in[4], zll_main_rotater1728_in[2], zll_main_rotater1728_in[1], zll_main_rotater1728_in[0]};
  assign zll_main_rotater1719_in = {zll_main_rotater17_in[31], zll_main_rotater17_in[30], zll_main_rotater17_in[29], zll_main_rotater17_in[28], zll_main_rotater17_in[27], zll_main_rotater17_in[26], zll_main_rotater17_in[25], zll_main_rotater17_in[24], zll_main_rotater17_in[23], zll_main_rotater17_in[22], zll_main_rotater17_in[21], zll_main_rotater17_in[20], zll_main_rotater17_in[19], zll_main_rotater17_in[18], zll_main_rotater17_in[17], zll_main_rotater17_in[16], zll_main_rotater17_in[15], zll_main_rotater17_in[14], zll_main_rotater17_in[13], zll_main_rotater17_in[12], zll_main_rotater17_in[11], zll_main_rotater17_in[10], zll_main_rotater17_in[9], zll_main_rotater17_in[8], zll_main_rotater17_in[7], zll_main_rotater17_in[6], zll_main_rotater17_in[5], zll_main_rotater17_in[2], zll_main_rotater17_in[4], zll_main_rotater17_in[3], zll_main_rotater17_in[1], zll_main_rotater17_in[0]};
  assign zll_main_rotater174_in = {zll_main_rotater1719_in[31], zll_main_rotater1719_in[30], zll_main_rotater1719_in[29], zll_main_rotater1719_in[28], zll_main_rotater1719_in[27], zll_main_rotater1719_in[26], zll_main_rotater1719_in[1], zll_main_rotater1719_in[25], zll_main_rotater1719_in[24], zll_main_rotater1719_in[23], zll_main_rotater1719_in[22], zll_main_rotater1719_in[21], zll_main_rotater1719_in[20], zll_main_rotater1719_in[19], zll_main_rotater1719_in[18], zll_main_rotater1719_in[17], zll_main_rotater1719_in[16], zll_main_rotater1719_in[15], zll_main_rotater1719_in[14], zll_main_rotater1719_in[13], zll_main_rotater1719_in[12], zll_main_rotater1719_in[11], zll_main_rotater1719_in[10], zll_main_rotater1719_in[9], zll_main_rotater1719_in[8], zll_main_rotater1719_in[7], zll_main_rotater1719_in[6], zll_main_rotater1719_in[5], zll_main_rotater1719_in[4], zll_main_rotater1719_in[3], zll_main_rotater1719_in[2], zll_main_rotater1719_in[0]};
  assign main_rotater19_in = main_sigma1_in[31:0];
  assign zll_main_rotater1931_in = main_rotater19_in[31:0];
  assign zll_main_rotater1912_in = {zll_main_rotater1931_in[30], zll_main_rotater1931_in[31], zll_main_rotater1931_in[29], zll_main_rotater1931_in[28], zll_main_rotater1931_in[27], zll_main_rotater1931_in[26], zll_main_rotater1931_in[25], zll_main_rotater1931_in[24], zll_main_rotater1931_in[23], zll_main_rotater1931_in[22], zll_main_rotater1931_in[21], zll_main_rotater1931_in[20], zll_main_rotater1931_in[19], zll_main_rotater1931_in[18], zll_main_rotater1931_in[17], zll_main_rotater1931_in[16], zll_main_rotater1931_in[15], zll_main_rotater1931_in[14], zll_main_rotater1931_in[13], zll_main_rotater1931_in[12], zll_main_rotater1931_in[11], zll_main_rotater1931_in[10], zll_main_rotater1931_in[9], zll_main_rotater1931_in[8], zll_main_rotater1931_in[7], zll_main_rotater1931_in[6], zll_main_rotater1931_in[5], zll_main_rotater1931_in[4], zll_main_rotater1931_in[3], zll_main_rotater1931_in[2], zll_main_rotater1931_in[1], zll_main_rotater1931_in[0]};
  assign zll_main_rotater198_in = {zll_main_rotater1912_in[27], zll_main_rotater1912_in[31], zll_main_rotater1912_in[30], zll_main_rotater1912_in[29], zll_main_rotater1912_in[28], zll_main_rotater1912_in[26], zll_main_rotater1912_in[25], zll_main_rotater1912_in[24], zll_main_rotater1912_in[23], zll_main_rotater1912_in[22], zll_main_rotater1912_in[21], zll_main_rotater1912_in[20], zll_main_rotater1912_in[19], zll_main_rotater1912_in[18], zll_main_rotater1912_in[17], zll_main_rotater1912_in[16], zll_main_rotater1912_in[15], zll_main_rotater1912_in[14], zll_main_rotater1912_in[13], zll_main_rotater1912_in[12], zll_main_rotater1912_in[11], zll_main_rotater1912_in[10], zll_main_rotater1912_in[9], zll_main_rotater1912_in[8], zll_main_rotater1912_in[7], zll_main_rotater1912_in[6], zll_main_rotater1912_in[5], zll_main_rotater1912_in[4], zll_main_rotater1912_in[3], zll_main_rotater1912_in[2], zll_main_rotater1912_in[1], zll_main_rotater1912_in[0]};
  assign zll_main_rotater1911_in = {zll_main_rotater198_in[26], zll_main_rotater198_in[31], zll_main_rotater198_in[30], zll_main_rotater198_in[29], zll_main_rotater198_in[28], zll_main_rotater198_in[27], zll_main_rotater198_in[25], zll_main_rotater198_in[24], zll_main_rotater198_in[23], zll_main_rotater198_in[22], zll_main_rotater198_in[21], zll_main_rotater198_in[20], zll_main_rotater198_in[19], zll_main_rotater198_in[18], zll_main_rotater198_in[17], zll_main_rotater198_in[16], zll_main_rotater198_in[15], zll_main_rotater198_in[14], zll_main_rotater198_in[13], zll_main_rotater198_in[12], zll_main_rotater198_in[11], zll_main_rotater198_in[10], zll_main_rotater198_in[9], zll_main_rotater198_in[8], zll_main_rotater198_in[7], zll_main_rotater198_in[6], zll_main_rotater198_in[5], zll_main_rotater198_in[4], zll_main_rotater198_in[3], zll_main_rotater198_in[2], zll_main_rotater198_in[1], zll_main_rotater198_in[0]};
  assign zll_main_rotater1929_in = {zll_main_rotater1911_in[31], zll_main_rotater1911_in[30], zll_main_rotater1911_in[29], zll_main_rotater1911_in[28], zll_main_rotater1911_in[24], zll_main_rotater1911_in[27], zll_main_rotater1911_in[26], zll_main_rotater1911_in[25], zll_main_rotater1911_in[23], zll_main_rotater1911_in[22], zll_main_rotater1911_in[21], zll_main_rotater1911_in[20], zll_main_rotater1911_in[19], zll_main_rotater1911_in[18], zll_main_rotater1911_in[17], zll_main_rotater1911_in[16], zll_main_rotater1911_in[15], zll_main_rotater1911_in[14], zll_main_rotater1911_in[13], zll_main_rotater1911_in[12], zll_main_rotater1911_in[11], zll_main_rotater1911_in[10], zll_main_rotater1911_in[9], zll_main_rotater1911_in[8], zll_main_rotater1911_in[7], zll_main_rotater1911_in[6], zll_main_rotater1911_in[5], zll_main_rotater1911_in[4], zll_main_rotater1911_in[3], zll_main_rotater1911_in[2], zll_main_rotater1911_in[1], zll_main_rotater1911_in[0]};
  assign zll_main_rotater194_in = {zll_main_rotater1929_in[31], zll_main_rotater1929_in[23], zll_main_rotater1929_in[30], zll_main_rotater1929_in[29], zll_main_rotater1929_in[28], zll_main_rotater1929_in[27], zll_main_rotater1929_in[26], zll_main_rotater1929_in[25], zll_main_rotater1929_in[24], zll_main_rotater1929_in[22], zll_main_rotater1929_in[21], zll_main_rotater1929_in[20], zll_main_rotater1929_in[19], zll_main_rotater1929_in[18], zll_main_rotater1929_in[17], zll_main_rotater1929_in[16], zll_main_rotater1929_in[15], zll_main_rotater1929_in[14], zll_main_rotater1929_in[13], zll_main_rotater1929_in[12], zll_main_rotater1929_in[11], zll_main_rotater1929_in[10], zll_main_rotater1929_in[9], zll_main_rotater1929_in[8], zll_main_rotater1929_in[7], zll_main_rotater1929_in[6], zll_main_rotater1929_in[5], zll_main_rotater1929_in[4], zll_main_rotater1929_in[3], zll_main_rotater1929_in[2], zll_main_rotater1929_in[1], zll_main_rotater1929_in[0]};
  assign zll_main_rotater1930_in = {zll_main_rotater194_in[31], zll_main_rotater194_in[30], zll_main_rotater194_in[29], zll_main_rotater194_in[28], zll_main_rotater194_in[27], zll_main_rotater194_in[26], zll_main_rotater194_in[25], zll_main_rotater194_in[24], zll_main_rotater194_in[22], zll_main_rotater194_in[23], zll_main_rotater194_in[21], zll_main_rotater194_in[20], zll_main_rotater194_in[19], zll_main_rotater194_in[18], zll_main_rotater194_in[17], zll_main_rotater194_in[16], zll_main_rotater194_in[15], zll_main_rotater194_in[14], zll_main_rotater194_in[13], zll_main_rotater194_in[12], zll_main_rotater194_in[11], zll_main_rotater194_in[10], zll_main_rotater194_in[9], zll_main_rotater194_in[8], zll_main_rotater194_in[7], zll_main_rotater194_in[6], zll_main_rotater194_in[5], zll_main_rotater194_in[4], zll_main_rotater194_in[3], zll_main_rotater194_in[2], zll_main_rotater194_in[1], zll_main_rotater194_in[0]};
  assign zll_main_rotater1918_in = {zll_main_rotater1930_in[31], zll_main_rotater1930_in[30], zll_main_rotater1930_in[29], zll_main_rotater1930_in[28], zll_main_rotater1930_in[27], zll_main_rotater1930_in[26], zll_main_rotater1930_in[25], zll_main_rotater1930_in[24], zll_main_rotater1930_in[23], zll_main_rotater1930_in[21], zll_main_rotater1930_in[22], zll_main_rotater1930_in[20], zll_main_rotater1930_in[19], zll_main_rotater1930_in[18], zll_main_rotater1930_in[17], zll_main_rotater1930_in[16], zll_main_rotater1930_in[15], zll_main_rotater1930_in[14], zll_main_rotater1930_in[13], zll_main_rotater1930_in[12], zll_main_rotater1930_in[11], zll_main_rotater1930_in[10], zll_main_rotater1930_in[9], zll_main_rotater1930_in[8], zll_main_rotater1930_in[7], zll_main_rotater1930_in[6], zll_main_rotater1930_in[5], zll_main_rotater1930_in[4], zll_main_rotater1930_in[3], zll_main_rotater1930_in[2], zll_main_rotater1930_in[1], zll_main_rotater1930_in[0]};
  assign zll_main_rotater1920_in = {zll_main_rotater1918_in[31], zll_main_rotater1918_in[30], zll_main_rotater1918_in[29], zll_main_rotater1918_in[28], zll_main_rotater1918_in[27], zll_main_rotater1918_in[26], zll_main_rotater1918_in[25], zll_main_rotater1918_in[24], zll_main_rotater1918_in[23], zll_main_rotater1918_in[22], zll_main_rotater1918_in[21], zll_main_rotater1918_in[19], zll_main_rotater1918_in[20], zll_main_rotater1918_in[18], zll_main_rotater1918_in[17], zll_main_rotater1918_in[16], zll_main_rotater1918_in[15], zll_main_rotater1918_in[14], zll_main_rotater1918_in[13], zll_main_rotater1918_in[12], zll_main_rotater1918_in[11], zll_main_rotater1918_in[10], zll_main_rotater1918_in[9], zll_main_rotater1918_in[8], zll_main_rotater1918_in[7], zll_main_rotater1918_in[6], zll_main_rotater1918_in[5], zll_main_rotater1918_in[4], zll_main_rotater1918_in[3], zll_main_rotater1918_in[2], zll_main_rotater1918_in[1], zll_main_rotater1918_in[0]};
  assign zll_main_rotater196_in = {zll_main_rotater1920_in[31], zll_main_rotater1920_in[30], zll_main_rotater1920_in[29], zll_main_rotater1920_in[28], zll_main_rotater1920_in[27], zll_main_rotater1920_in[17], zll_main_rotater1920_in[26], zll_main_rotater1920_in[25], zll_main_rotater1920_in[24], zll_main_rotater1920_in[23], zll_main_rotater1920_in[22], zll_main_rotater1920_in[21], zll_main_rotater1920_in[20], zll_main_rotater1920_in[19], zll_main_rotater1920_in[18], zll_main_rotater1920_in[16], zll_main_rotater1920_in[15], zll_main_rotater1920_in[14], zll_main_rotater1920_in[13], zll_main_rotater1920_in[12], zll_main_rotater1920_in[11], zll_main_rotater1920_in[10], zll_main_rotater1920_in[9], zll_main_rotater1920_in[8], zll_main_rotater1920_in[7], zll_main_rotater1920_in[6], zll_main_rotater1920_in[5], zll_main_rotater1920_in[4], zll_main_rotater1920_in[3], zll_main_rotater1920_in[2], zll_main_rotater1920_in[1], zll_main_rotater1920_in[0]};
  assign zll_main_rotater1924_in = {zll_main_rotater196_in[31], zll_main_rotater196_in[30], zll_main_rotater196_in[29], zll_main_rotater196_in[28], zll_main_rotater196_in[27], zll_main_rotater196_in[16], zll_main_rotater196_in[26], zll_main_rotater196_in[25], zll_main_rotater196_in[24], zll_main_rotater196_in[23], zll_main_rotater196_in[22], zll_main_rotater196_in[21], zll_main_rotater196_in[20], zll_main_rotater196_in[19], zll_main_rotater196_in[18], zll_main_rotater196_in[17], zll_main_rotater196_in[15], zll_main_rotater196_in[14], zll_main_rotater196_in[13], zll_main_rotater196_in[12], zll_main_rotater196_in[11], zll_main_rotater196_in[10], zll_main_rotater196_in[9], zll_main_rotater196_in[8], zll_main_rotater196_in[7], zll_main_rotater196_in[6], zll_main_rotater196_in[5], zll_main_rotater196_in[4], zll_main_rotater196_in[3], zll_main_rotater196_in[2], zll_main_rotater196_in[1], zll_main_rotater196_in[0]};
  assign zll_main_rotater1923_in = {zll_main_rotater1924_in[31], zll_main_rotater1924_in[30], zll_main_rotater1924_in[29], zll_main_rotater1924_in[28], zll_main_rotater1924_in[27], zll_main_rotater1924_in[15], zll_main_rotater1924_in[26], zll_main_rotater1924_in[25], zll_main_rotater1924_in[24], zll_main_rotater1924_in[23], zll_main_rotater1924_in[22], zll_main_rotater1924_in[21], zll_main_rotater1924_in[20], zll_main_rotater1924_in[19], zll_main_rotater1924_in[18], zll_main_rotater1924_in[17], zll_main_rotater1924_in[16], zll_main_rotater1924_in[14], zll_main_rotater1924_in[13], zll_main_rotater1924_in[12], zll_main_rotater1924_in[11], zll_main_rotater1924_in[10], zll_main_rotater1924_in[9], zll_main_rotater1924_in[8], zll_main_rotater1924_in[7], zll_main_rotater1924_in[6], zll_main_rotater1924_in[5], zll_main_rotater1924_in[4], zll_main_rotater1924_in[3], zll_main_rotater1924_in[2], zll_main_rotater1924_in[1], zll_main_rotater1924_in[0]};
  assign zll_main_rotater1916_in = {zll_main_rotater1923_in[31], zll_main_rotater1923_in[30], zll_main_rotater1923_in[29], zll_main_rotater1923_in[28], zll_main_rotater1923_in[27], zll_main_rotater1923_in[26], zll_main_rotater1923_in[25], zll_main_rotater1923_in[24], zll_main_rotater1923_in[23], zll_main_rotater1923_in[22], zll_main_rotater1923_in[21], zll_main_rotater1923_in[20], zll_main_rotater1923_in[19], zll_main_rotater1923_in[18], zll_main_rotater1923_in[17], zll_main_rotater1923_in[14], zll_main_rotater1923_in[16], zll_main_rotater1923_in[15], zll_main_rotater1923_in[13], zll_main_rotater1923_in[12], zll_main_rotater1923_in[11], zll_main_rotater1923_in[10], zll_main_rotater1923_in[9], zll_main_rotater1923_in[8], zll_main_rotater1923_in[7], zll_main_rotater1923_in[6], zll_main_rotater1923_in[5], zll_main_rotater1923_in[4], zll_main_rotater1923_in[3], zll_main_rotater1923_in[2], zll_main_rotater1923_in[1], zll_main_rotater1923_in[0]};
  assign zll_main_rotater1919_in = {zll_main_rotater1916_in[31], zll_main_rotater1916_in[30], zll_main_rotater1916_in[29], zll_main_rotater1916_in[28], zll_main_rotater1916_in[27], zll_main_rotater1916_in[26], zll_main_rotater1916_in[25], zll_main_rotater1916_in[24], zll_main_rotater1916_in[23], zll_main_rotater1916_in[22], zll_main_rotater1916_in[21], zll_main_rotater1916_in[20], zll_main_rotater1916_in[13], zll_main_rotater1916_in[19], zll_main_rotater1916_in[18], zll_main_rotater1916_in[17], zll_main_rotater1916_in[16], zll_main_rotater1916_in[15], zll_main_rotater1916_in[14], zll_main_rotater1916_in[12], zll_main_rotater1916_in[11], zll_main_rotater1916_in[10], zll_main_rotater1916_in[9], zll_main_rotater1916_in[8], zll_main_rotater1916_in[7], zll_main_rotater1916_in[6], zll_main_rotater1916_in[5], zll_main_rotater1916_in[4], zll_main_rotater1916_in[3], zll_main_rotater1916_in[2], zll_main_rotater1916_in[1], zll_main_rotater1916_in[0]};
  assign zll_main_rotater1917_in = {zll_main_rotater1919_in[31], zll_main_rotater1919_in[30], zll_main_rotater1919_in[29], zll_main_rotater1919_in[28], zll_main_rotater1919_in[27], zll_main_rotater1919_in[26], zll_main_rotater1919_in[25], zll_main_rotater1919_in[24], zll_main_rotater1919_in[23], zll_main_rotater1919_in[22], zll_main_rotater1919_in[21], zll_main_rotater1919_in[20], zll_main_rotater1919_in[19], zll_main_rotater1919_in[18], zll_main_rotater1919_in[17], zll_main_rotater1919_in[16], zll_main_rotater1919_in[12], zll_main_rotater1919_in[15], zll_main_rotater1919_in[14], zll_main_rotater1919_in[13], zll_main_rotater1919_in[11], zll_main_rotater1919_in[10], zll_main_rotater1919_in[9], zll_main_rotater1919_in[8], zll_main_rotater1919_in[7], zll_main_rotater1919_in[6], zll_main_rotater1919_in[5], zll_main_rotater1919_in[4], zll_main_rotater1919_in[3], zll_main_rotater1919_in[2], zll_main_rotater1919_in[1], zll_main_rotater1919_in[0]};
  assign zll_main_rotater1926_in = {zll_main_rotater1917_in[11], zll_main_rotater1917_in[31], zll_main_rotater1917_in[30], zll_main_rotater1917_in[29], zll_main_rotater1917_in[28], zll_main_rotater1917_in[27], zll_main_rotater1917_in[26], zll_main_rotater1917_in[25], zll_main_rotater1917_in[24], zll_main_rotater1917_in[23], zll_main_rotater1917_in[22], zll_main_rotater1917_in[21], zll_main_rotater1917_in[20], zll_main_rotater1917_in[19], zll_main_rotater1917_in[18], zll_main_rotater1917_in[17], zll_main_rotater1917_in[16], zll_main_rotater1917_in[15], zll_main_rotater1917_in[14], zll_main_rotater1917_in[13], zll_main_rotater1917_in[12], zll_main_rotater1917_in[10], zll_main_rotater1917_in[9], zll_main_rotater1917_in[8], zll_main_rotater1917_in[7], zll_main_rotater1917_in[6], zll_main_rotater1917_in[5], zll_main_rotater1917_in[4], zll_main_rotater1917_in[3], zll_main_rotater1917_in[2], zll_main_rotater1917_in[1], zll_main_rotater1917_in[0]};
  assign zll_main_rotater195_in = {zll_main_rotater1926_in[31], zll_main_rotater1926_in[30], zll_main_rotater1926_in[29], zll_main_rotater1926_in[10], zll_main_rotater1926_in[28], zll_main_rotater1926_in[27], zll_main_rotater1926_in[26], zll_main_rotater1926_in[25], zll_main_rotater1926_in[24], zll_main_rotater1926_in[23], zll_main_rotater1926_in[22], zll_main_rotater1926_in[21], zll_main_rotater1926_in[20], zll_main_rotater1926_in[19], zll_main_rotater1926_in[18], zll_main_rotater1926_in[17], zll_main_rotater1926_in[16], zll_main_rotater1926_in[15], zll_main_rotater1926_in[14], zll_main_rotater1926_in[13], zll_main_rotater1926_in[12], zll_main_rotater1926_in[11], zll_main_rotater1926_in[9], zll_main_rotater1926_in[8], zll_main_rotater1926_in[7], zll_main_rotater1926_in[6], zll_main_rotater1926_in[5], zll_main_rotater1926_in[4], zll_main_rotater1926_in[3], zll_main_rotater1926_in[2], zll_main_rotater1926_in[1], zll_main_rotater1926_in[0]};
  assign zll_main_rotater1914_in = {zll_main_rotater195_in[9], zll_main_rotater195_in[31], zll_main_rotater195_in[30], zll_main_rotater195_in[29], zll_main_rotater195_in[28], zll_main_rotater195_in[27], zll_main_rotater195_in[26], zll_main_rotater195_in[25], zll_main_rotater195_in[24], zll_main_rotater195_in[23], zll_main_rotater195_in[22], zll_main_rotater195_in[21], zll_main_rotater195_in[20], zll_main_rotater195_in[19], zll_main_rotater195_in[18], zll_main_rotater195_in[17], zll_main_rotater195_in[16], zll_main_rotater195_in[15], zll_main_rotater195_in[14], zll_main_rotater195_in[13], zll_main_rotater195_in[12], zll_main_rotater195_in[11], zll_main_rotater195_in[10], zll_main_rotater195_in[8], zll_main_rotater195_in[7], zll_main_rotater195_in[6], zll_main_rotater195_in[5], zll_main_rotater195_in[4], zll_main_rotater195_in[3], zll_main_rotater195_in[2], zll_main_rotater195_in[1], zll_main_rotater195_in[0]};
  assign zll_main_rotater193_in = {zll_main_rotater1914_in[31], zll_main_rotater1914_in[30], zll_main_rotater1914_in[29], zll_main_rotater1914_in[28], zll_main_rotater1914_in[27], zll_main_rotater1914_in[26], zll_main_rotater1914_in[25], zll_main_rotater1914_in[24], zll_main_rotater1914_in[23], zll_main_rotater1914_in[22], zll_main_rotater1914_in[21], zll_main_rotater1914_in[20], zll_main_rotater1914_in[19], zll_main_rotater1914_in[18], zll_main_rotater1914_in[17], zll_main_rotater1914_in[16], zll_main_rotater1914_in[15], zll_main_rotater1914_in[14], zll_main_rotater1914_in[13], zll_main_rotater1914_in[12], zll_main_rotater1914_in[8], zll_main_rotater1914_in[11], zll_main_rotater1914_in[10], zll_main_rotater1914_in[9], zll_main_rotater1914_in[7], zll_main_rotater1914_in[6], zll_main_rotater1914_in[5], zll_main_rotater1914_in[4], zll_main_rotater1914_in[3], zll_main_rotater1914_in[2], zll_main_rotater1914_in[1], zll_main_rotater1914_in[0]};
  assign zll_main_rotater192_in = {zll_main_rotater193_in[7], zll_main_rotater193_in[31], zll_main_rotater193_in[30], zll_main_rotater193_in[29], zll_main_rotater193_in[28], zll_main_rotater193_in[27], zll_main_rotater193_in[26], zll_main_rotater193_in[25], zll_main_rotater193_in[24], zll_main_rotater193_in[23], zll_main_rotater193_in[22], zll_main_rotater193_in[21], zll_main_rotater193_in[20], zll_main_rotater193_in[19], zll_main_rotater193_in[18], zll_main_rotater193_in[17], zll_main_rotater193_in[16], zll_main_rotater193_in[15], zll_main_rotater193_in[14], zll_main_rotater193_in[13], zll_main_rotater193_in[12], zll_main_rotater193_in[11], zll_main_rotater193_in[10], zll_main_rotater193_in[9], zll_main_rotater193_in[8], zll_main_rotater193_in[6], zll_main_rotater193_in[5], zll_main_rotater193_in[4], zll_main_rotater193_in[3], zll_main_rotater193_in[2], zll_main_rotater193_in[1], zll_main_rotater193_in[0]};
  assign zll_main_rotater197_in = {zll_main_rotater192_in[31], zll_main_rotater192_in[30], zll_main_rotater192_in[29], zll_main_rotater192_in[28], zll_main_rotater192_in[27], zll_main_rotater192_in[26], zll_main_rotater192_in[25], zll_main_rotater192_in[24], zll_main_rotater192_in[23], zll_main_rotater192_in[22], zll_main_rotater192_in[21], zll_main_rotater192_in[20], zll_main_rotater192_in[19], zll_main_rotater192_in[18], zll_main_rotater192_in[17], zll_main_rotater192_in[16], zll_main_rotater192_in[15], zll_main_rotater192_in[14], zll_main_rotater192_in[13], zll_main_rotater192_in[12], zll_main_rotater192_in[5], zll_main_rotater192_in[11], zll_main_rotater192_in[10], zll_main_rotater192_in[9], zll_main_rotater192_in[8], zll_main_rotater192_in[7], zll_main_rotater192_in[6], zll_main_rotater192_in[4], zll_main_rotater192_in[3], zll_main_rotater192_in[2], zll_main_rotater192_in[1], zll_main_rotater192_in[0]};
  assign zll_main_rotater19_in = {zll_main_rotater197_in[31], zll_main_rotater197_in[4], zll_main_rotater197_in[30], zll_main_rotater197_in[29], zll_main_rotater197_in[28], zll_main_rotater197_in[27], zll_main_rotater197_in[26], zll_main_rotater197_in[25], zll_main_rotater197_in[24], zll_main_rotater197_in[23], zll_main_rotater197_in[22], zll_main_rotater197_in[21], zll_main_rotater197_in[20], zll_main_rotater197_in[19], zll_main_rotater197_in[18], zll_main_rotater197_in[17], zll_main_rotater197_in[16], zll_main_rotater197_in[15], zll_main_rotater197_in[14], zll_main_rotater197_in[13], zll_main_rotater197_in[12], zll_main_rotater197_in[11], zll_main_rotater197_in[10], zll_main_rotater197_in[9], zll_main_rotater197_in[8], zll_main_rotater197_in[7], zll_main_rotater197_in[6], zll_main_rotater197_in[5], zll_main_rotater197_in[3], zll_main_rotater197_in[2], zll_main_rotater197_in[1], zll_main_rotater197_in[0]};
  assign zll_main_rotater199_in = {zll_main_rotater19_in[31], zll_main_rotater19_in[30], zll_main_rotater19_in[29], zll_main_rotater19_in[28], zll_main_rotater19_in[27], zll_main_rotater19_in[26], zll_main_rotater19_in[25], zll_main_rotater19_in[24], zll_main_rotater19_in[23], zll_main_rotater19_in[3], zll_main_rotater19_in[22], zll_main_rotater19_in[21], zll_main_rotater19_in[20], zll_main_rotater19_in[19], zll_main_rotater19_in[18], zll_main_rotater19_in[17], zll_main_rotater19_in[16], zll_main_rotater19_in[15], zll_main_rotater19_in[14], zll_main_rotater19_in[13], zll_main_rotater19_in[12], zll_main_rotater19_in[11], zll_main_rotater19_in[10], zll_main_rotater19_in[9], zll_main_rotater19_in[8], zll_main_rotater19_in[7], zll_main_rotater19_in[6], zll_main_rotater19_in[5], zll_main_rotater19_in[4], zll_main_rotater19_in[2], zll_main_rotater19_in[1], zll_main_rotater19_in[0]};
  assign zll_main_rotater1928_in = {zll_main_rotater199_in[31], zll_main_rotater199_in[30], zll_main_rotater199_in[29], zll_main_rotater199_in[28], zll_main_rotater199_in[27], zll_main_rotater199_in[26], zll_main_rotater199_in[25], zll_main_rotater199_in[24], zll_main_rotater199_in[23], zll_main_rotater199_in[22], zll_main_rotater199_in[21], zll_main_rotater199_in[20], zll_main_rotater199_in[19], zll_main_rotater199_in[18], zll_main_rotater199_in[17], zll_main_rotater199_in[16], zll_main_rotater199_in[15], zll_main_rotater199_in[14], zll_main_rotater199_in[13], zll_main_rotater199_in[2], zll_main_rotater199_in[12], zll_main_rotater199_in[11], zll_main_rotater199_in[10], zll_main_rotater199_in[9], zll_main_rotater199_in[8], zll_main_rotater199_in[7], zll_main_rotater199_in[6], zll_main_rotater199_in[5], zll_main_rotater199_in[4], zll_main_rotater199_in[3], zll_main_rotater199_in[1], zll_main_rotater199_in[0]};
  assign zll_main_rotater1910_in = {zll_main_rotater1928_in[31], zll_main_rotater1928_in[30], zll_main_rotater1928_in[29], zll_main_rotater1928_in[28], zll_main_rotater1928_in[27], zll_main_rotater1928_in[26], zll_main_rotater1928_in[25], zll_main_rotater1928_in[24], zll_main_rotater1928_in[23], zll_main_rotater1928_in[22], zll_main_rotater1928_in[21], zll_main_rotater1928_in[20], zll_main_rotater1928_in[19], zll_main_rotater1928_in[18], zll_main_rotater1928_in[17], zll_main_rotater1928_in[16], zll_main_rotater1928_in[15], zll_main_rotater1928_in[14], zll_main_rotater1928_in[13], zll_main_rotater1928_in[12], zll_main_rotater1928_in[11], zll_main_rotater1928_in[10], zll_main_rotater1928_in[9], zll_main_rotater1928_in[8], zll_main_rotater1928_in[7], zll_main_rotater1928_in[6], zll_main_rotater1928_in[5], zll_main_rotater1928_in[1], zll_main_rotater1928_in[4], zll_main_rotater1928_in[3], zll_main_rotater1928_in[2], zll_main_rotater1928_in[0]};
  assign xorw32_in = {{zll_main_rotater174_in[8], zll_main_rotater174_in[15], zll_main_rotater174_in[27], zll_main_rotater174_in[5], zll_main_rotater174_in[1], zll_main_rotater174_in[14], zll_main_rotater174_in[9], zll_main_rotater174_in[10], zll_main_rotater174_in[26], zll_main_rotater174_in[7], zll_main_rotater174_in[17], zll_main_rotater174_in[13], zll_main_rotater174_in[22], zll_main_rotater174_in[30], zll_main_rotater174_in[3], zll_main_rotater174_in[25], zll_main_rotater174_in[0], zll_main_rotater174_in[31], zll_main_rotater174_in[16], zll_main_rotater174_in[19], zll_main_rotater174_in[29], zll_main_rotater174_in[24], zll_main_rotater174_in[20], zll_main_rotater174_in[6], zll_main_rotater174_in[11], zll_main_rotater174_in[4], zll_main_rotater174_in[21], zll_main_rotater174_in[18], zll_main_rotater174_in[28], zll_main_rotater174_in[2], zll_main_rotater174_in[23], zll_main_rotater174_in[12]}, {zll_main_rotater1910_in[2], zll_main_rotater1910_in[18], zll_main_rotater1910_in[19], zll_main_rotater1910_in[20], zll_main_rotater1910_in[5], zll_main_rotater1910_in[13], zll_main_rotater1910_in[7], zll_main_rotater1910_in[28], zll_main_rotater1910_in[25], zll_main_rotater1910_in[29], zll_main_rotater1910_in[6], zll_main_rotater1910_in[31], zll_main_rotater1910_in[1], zll_main_rotater1910_in[8], zll_main_rotater1910_in[30], zll_main_rotater1910_in[22], zll_main_rotater1910_in[12], zll_main_rotater1910_in[4], zll_main_rotater1910_in[0], zll_main_rotater1910_in[21], zll_main_rotater1910_in[23], zll_main_rotater1910_in[16], zll_main_rotater1910_in[15], zll_main_rotater1910_in[24], zll_main_rotater1910_in[27], zll_main_rotater1910_in[10], zll_main_rotater1910_in[17], zll_main_rotater1910_in[26], zll_main_rotater1910_in[14], zll_main_rotater1910_in[11], zll_main_rotater1910_in[3], zll_main_rotater1910_in[9]}};
  xorW32  inst (xorw32_in[63:32], xorw32_in[31:0], extres[31:0]);
  assign main_shiftr10_in = main_sigma1_in[31:0];
  assign zll_main_shiftr1028_in = main_shiftr10_in[31:0];
  assign zll_main_shiftr109_in = {zll_main_shiftr1028_in[29], zll_main_shiftr1028_in[31], zll_main_shiftr1028_in[30], zll_main_shiftr1028_in[28], zll_main_shiftr1028_in[27], zll_main_shiftr1028_in[26], zll_main_shiftr1028_in[25], zll_main_shiftr1028_in[24], zll_main_shiftr1028_in[23], zll_main_shiftr1028_in[22], zll_main_shiftr1028_in[21], zll_main_shiftr1028_in[20], zll_main_shiftr1028_in[19], zll_main_shiftr1028_in[18], zll_main_shiftr1028_in[17], zll_main_shiftr1028_in[16], zll_main_shiftr1028_in[15], zll_main_shiftr1028_in[14], zll_main_shiftr1028_in[13], zll_main_shiftr1028_in[12], zll_main_shiftr1028_in[11], zll_main_shiftr1028_in[10], zll_main_shiftr1028_in[9], zll_main_shiftr1028_in[8], zll_main_shiftr1028_in[7], zll_main_shiftr1028_in[6], zll_main_shiftr1028_in[5], zll_main_shiftr1028_in[4], zll_main_shiftr1028_in[3], zll_main_shiftr1028_in[2], zll_main_shiftr1028_in[1], zll_main_shiftr1028_in[0]};
  assign zll_main_shiftr105_in = {zll_main_shiftr109_in[31], zll_main_shiftr109_in[30], zll_main_shiftr109_in[29], zll_main_shiftr109_in[27], zll_main_shiftr109_in[28], zll_main_shiftr109_in[26], zll_main_shiftr109_in[25], zll_main_shiftr109_in[24], zll_main_shiftr109_in[23], zll_main_shiftr109_in[22], zll_main_shiftr109_in[21], zll_main_shiftr109_in[20], zll_main_shiftr109_in[19], zll_main_shiftr109_in[18], zll_main_shiftr109_in[17], zll_main_shiftr109_in[16], zll_main_shiftr109_in[15], zll_main_shiftr109_in[14], zll_main_shiftr109_in[13], zll_main_shiftr109_in[12], zll_main_shiftr109_in[11], zll_main_shiftr109_in[10], zll_main_shiftr109_in[9], zll_main_shiftr109_in[8], zll_main_shiftr109_in[7], zll_main_shiftr109_in[6], zll_main_shiftr109_in[5], zll_main_shiftr109_in[4], zll_main_shiftr109_in[3], zll_main_shiftr109_in[2], zll_main_shiftr109_in[1], zll_main_shiftr109_in[0]};
  assign zll_main_shiftr10_in = {zll_main_shiftr105_in[31], zll_main_shiftr105_in[26], zll_main_shiftr105_in[30], zll_main_shiftr105_in[29], zll_main_shiftr105_in[28], zll_main_shiftr105_in[27], zll_main_shiftr105_in[25], zll_main_shiftr105_in[24], zll_main_shiftr105_in[23], zll_main_shiftr105_in[22], zll_main_shiftr105_in[21], zll_main_shiftr105_in[20], zll_main_shiftr105_in[19], zll_main_shiftr105_in[18], zll_main_shiftr105_in[17], zll_main_shiftr105_in[16], zll_main_shiftr105_in[15], zll_main_shiftr105_in[14], zll_main_shiftr105_in[13], zll_main_shiftr105_in[12], zll_main_shiftr105_in[11], zll_main_shiftr105_in[10], zll_main_shiftr105_in[9], zll_main_shiftr105_in[8], zll_main_shiftr105_in[7], zll_main_shiftr105_in[6], zll_main_shiftr105_in[5], zll_main_shiftr105_in[4], zll_main_shiftr105_in[3], zll_main_shiftr105_in[2], zll_main_shiftr105_in[1], zll_main_shiftr105_in[0]};
  assign zll_main_shiftr1013_in = {zll_main_shiftr10_in[31], zll_main_shiftr10_in[30], zll_main_shiftr10_in[29], zll_main_shiftr10_in[24], zll_main_shiftr10_in[28], zll_main_shiftr10_in[27], zll_main_shiftr10_in[26], zll_main_shiftr10_in[25], zll_main_shiftr10_in[23], zll_main_shiftr10_in[22], zll_main_shiftr10_in[21], zll_main_shiftr10_in[20], zll_main_shiftr10_in[19], zll_main_shiftr10_in[18], zll_main_shiftr10_in[17], zll_main_shiftr10_in[16], zll_main_shiftr10_in[15], zll_main_shiftr10_in[14], zll_main_shiftr10_in[13], zll_main_shiftr10_in[12], zll_main_shiftr10_in[11], zll_main_shiftr10_in[10], zll_main_shiftr10_in[9], zll_main_shiftr10_in[8], zll_main_shiftr10_in[7], zll_main_shiftr10_in[6], zll_main_shiftr10_in[5], zll_main_shiftr10_in[4], zll_main_shiftr10_in[3], zll_main_shiftr10_in[2], zll_main_shiftr10_in[1], zll_main_shiftr10_in[0]};
  assign zll_main_shiftr108_in = {zll_main_shiftr1013_in[31], zll_main_shiftr1013_in[30], zll_main_shiftr1013_in[29], zll_main_shiftr1013_in[28], zll_main_shiftr1013_in[27], zll_main_shiftr1013_in[26], zll_main_shiftr1013_in[25], zll_main_shiftr1013_in[22], zll_main_shiftr1013_in[24], zll_main_shiftr1013_in[23], zll_main_shiftr1013_in[21], zll_main_shiftr1013_in[20], zll_main_shiftr1013_in[19], zll_main_shiftr1013_in[18], zll_main_shiftr1013_in[17], zll_main_shiftr1013_in[16], zll_main_shiftr1013_in[15], zll_main_shiftr1013_in[14], zll_main_shiftr1013_in[13], zll_main_shiftr1013_in[12], zll_main_shiftr1013_in[11], zll_main_shiftr1013_in[10], zll_main_shiftr1013_in[9], zll_main_shiftr1013_in[8], zll_main_shiftr1013_in[7], zll_main_shiftr1013_in[6], zll_main_shiftr1013_in[5], zll_main_shiftr1013_in[4], zll_main_shiftr1013_in[3], zll_main_shiftr1013_in[2], zll_main_shiftr1013_in[1], zll_main_shiftr1013_in[0]};
  assign zll_main_shiftr1011_in = {zll_main_shiftr108_in[31], zll_main_shiftr108_in[30], zll_main_shiftr108_in[29], zll_main_shiftr108_in[28], zll_main_shiftr108_in[27], zll_main_shiftr108_in[21], zll_main_shiftr108_in[26], zll_main_shiftr108_in[25], zll_main_shiftr108_in[24], zll_main_shiftr108_in[23], zll_main_shiftr108_in[22], zll_main_shiftr108_in[20], zll_main_shiftr108_in[19], zll_main_shiftr108_in[18], zll_main_shiftr108_in[17], zll_main_shiftr108_in[16], zll_main_shiftr108_in[15], zll_main_shiftr108_in[14], zll_main_shiftr108_in[13], zll_main_shiftr108_in[12], zll_main_shiftr108_in[11], zll_main_shiftr108_in[10], zll_main_shiftr108_in[9], zll_main_shiftr108_in[8], zll_main_shiftr108_in[7], zll_main_shiftr108_in[6], zll_main_shiftr108_in[5], zll_main_shiftr108_in[4], zll_main_shiftr108_in[3], zll_main_shiftr108_in[2], zll_main_shiftr108_in[1], zll_main_shiftr108_in[0]};
  assign zll_main_shiftr1016_in = {zll_main_shiftr1011_in[31], zll_main_shiftr1011_in[30], zll_main_shiftr1011_in[29], zll_main_shiftr1011_in[28], zll_main_shiftr1011_in[27], zll_main_shiftr1011_in[26], zll_main_shiftr1011_in[25], zll_main_shiftr1011_in[24], zll_main_shiftr1011_in[23], zll_main_shiftr1011_in[20], zll_main_shiftr1011_in[22], zll_main_shiftr1011_in[21], zll_main_shiftr1011_in[19], zll_main_shiftr1011_in[18], zll_main_shiftr1011_in[17], zll_main_shiftr1011_in[16], zll_main_shiftr1011_in[15], zll_main_shiftr1011_in[14], zll_main_shiftr1011_in[13], zll_main_shiftr1011_in[12], zll_main_shiftr1011_in[11], zll_main_shiftr1011_in[10], zll_main_shiftr1011_in[9], zll_main_shiftr1011_in[8], zll_main_shiftr1011_in[7], zll_main_shiftr1011_in[6], zll_main_shiftr1011_in[5], zll_main_shiftr1011_in[4], zll_main_shiftr1011_in[3], zll_main_shiftr1011_in[2], zll_main_shiftr1011_in[1], zll_main_shiftr1011_in[0]};
  assign zll_main_shiftr1021_in = {zll_main_shiftr1016_in[31], zll_main_shiftr1016_in[30], zll_main_shiftr1016_in[29], zll_main_shiftr1016_in[28], zll_main_shiftr1016_in[27], zll_main_shiftr1016_in[26], zll_main_shiftr1016_in[25], zll_main_shiftr1016_in[24], zll_main_shiftr1016_in[19], zll_main_shiftr1016_in[23], zll_main_shiftr1016_in[22], zll_main_shiftr1016_in[21], zll_main_shiftr1016_in[20], zll_main_shiftr1016_in[18], zll_main_shiftr1016_in[17], zll_main_shiftr1016_in[16], zll_main_shiftr1016_in[15], zll_main_shiftr1016_in[14], zll_main_shiftr1016_in[13], zll_main_shiftr1016_in[12], zll_main_shiftr1016_in[11], zll_main_shiftr1016_in[10], zll_main_shiftr1016_in[9], zll_main_shiftr1016_in[8], zll_main_shiftr1016_in[7], zll_main_shiftr1016_in[6], zll_main_shiftr1016_in[5], zll_main_shiftr1016_in[4], zll_main_shiftr1016_in[3], zll_main_shiftr1016_in[2], zll_main_shiftr1016_in[1], zll_main_shiftr1016_in[0]};
  assign zll_main_shiftr1024_in = {zll_main_shiftr1021_in[18], zll_main_shiftr1021_in[31], zll_main_shiftr1021_in[30], zll_main_shiftr1021_in[29], zll_main_shiftr1021_in[28], zll_main_shiftr1021_in[27], zll_main_shiftr1021_in[26], zll_main_shiftr1021_in[25], zll_main_shiftr1021_in[24], zll_main_shiftr1021_in[23], zll_main_shiftr1021_in[22], zll_main_shiftr1021_in[21], zll_main_shiftr1021_in[20], zll_main_shiftr1021_in[19], zll_main_shiftr1021_in[17], zll_main_shiftr1021_in[16], zll_main_shiftr1021_in[15], zll_main_shiftr1021_in[14], zll_main_shiftr1021_in[13], zll_main_shiftr1021_in[12], zll_main_shiftr1021_in[11], zll_main_shiftr1021_in[10], zll_main_shiftr1021_in[9], zll_main_shiftr1021_in[8], zll_main_shiftr1021_in[7], zll_main_shiftr1021_in[6], zll_main_shiftr1021_in[5], zll_main_shiftr1021_in[4], zll_main_shiftr1021_in[3], zll_main_shiftr1021_in[2], zll_main_shiftr1021_in[1], zll_main_shiftr1021_in[0]};
  assign zll_main_shiftr103_in = {zll_main_shiftr1024_in[31], zll_main_shiftr1024_in[30], zll_main_shiftr1024_in[29], zll_main_shiftr1024_in[28], zll_main_shiftr1024_in[27], zll_main_shiftr1024_in[26], zll_main_shiftr1024_in[25], zll_main_shiftr1024_in[24], zll_main_shiftr1024_in[23], zll_main_shiftr1024_in[22], zll_main_shiftr1024_in[21], zll_main_shiftr1024_in[20], zll_main_shiftr1024_in[19], zll_main_shiftr1024_in[17], zll_main_shiftr1024_in[18], zll_main_shiftr1024_in[16], zll_main_shiftr1024_in[15], zll_main_shiftr1024_in[14], zll_main_shiftr1024_in[13], zll_main_shiftr1024_in[12], zll_main_shiftr1024_in[11], zll_main_shiftr1024_in[10], zll_main_shiftr1024_in[9], zll_main_shiftr1024_in[8], zll_main_shiftr1024_in[7], zll_main_shiftr1024_in[6], zll_main_shiftr1024_in[5], zll_main_shiftr1024_in[4], zll_main_shiftr1024_in[3], zll_main_shiftr1024_in[2], zll_main_shiftr1024_in[1], zll_main_shiftr1024_in[0]};
  assign zll_main_shiftr106_in = {zll_main_shiftr103_in[31], zll_main_shiftr103_in[30], zll_main_shiftr103_in[29], zll_main_shiftr103_in[28], zll_main_shiftr103_in[27], zll_main_shiftr103_in[26], zll_main_shiftr103_in[25], zll_main_shiftr103_in[24], zll_main_shiftr103_in[23], zll_main_shiftr103_in[22], zll_main_shiftr103_in[16], zll_main_shiftr103_in[21], zll_main_shiftr103_in[20], zll_main_shiftr103_in[19], zll_main_shiftr103_in[18], zll_main_shiftr103_in[17], zll_main_shiftr103_in[15], zll_main_shiftr103_in[14], zll_main_shiftr103_in[13], zll_main_shiftr103_in[12], zll_main_shiftr103_in[11], zll_main_shiftr103_in[10], zll_main_shiftr103_in[9], zll_main_shiftr103_in[8], zll_main_shiftr103_in[7], zll_main_shiftr103_in[6], zll_main_shiftr103_in[5], zll_main_shiftr103_in[4], zll_main_shiftr103_in[3], zll_main_shiftr103_in[2], zll_main_shiftr103_in[1], zll_main_shiftr103_in[0]};
  assign zll_main_shiftr1017_in = {zll_main_shiftr106_in[31], zll_main_shiftr106_in[30], zll_main_shiftr106_in[29], zll_main_shiftr106_in[28], zll_main_shiftr106_in[27], zll_main_shiftr106_in[26], zll_main_shiftr106_in[15], zll_main_shiftr106_in[25], zll_main_shiftr106_in[24], zll_main_shiftr106_in[23], zll_main_shiftr106_in[22], zll_main_shiftr106_in[21], zll_main_shiftr106_in[20], zll_main_shiftr106_in[19], zll_main_shiftr106_in[18], zll_main_shiftr106_in[17], zll_main_shiftr106_in[16], zll_main_shiftr106_in[14], zll_main_shiftr106_in[13], zll_main_shiftr106_in[12], zll_main_shiftr106_in[11], zll_main_shiftr106_in[10], zll_main_shiftr106_in[9], zll_main_shiftr106_in[8], zll_main_shiftr106_in[7], zll_main_shiftr106_in[6], zll_main_shiftr106_in[5], zll_main_shiftr106_in[4], zll_main_shiftr106_in[3], zll_main_shiftr106_in[2], zll_main_shiftr106_in[1], zll_main_shiftr106_in[0]};
  assign zll_main_shiftr1012_in = {zll_main_shiftr1017_in[31], zll_main_shiftr1017_in[30], zll_main_shiftr1017_in[29], zll_main_shiftr1017_in[28], zll_main_shiftr1017_in[27], zll_main_shiftr1017_in[14], zll_main_shiftr1017_in[26], zll_main_shiftr1017_in[25], zll_main_shiftr1017_in[24], zll_main_shiftr1017_in[23], zll_main_shiftr1017_in[22], zll_main_shiftr1017_in[21], zll_main_shiftr1017_in[20], zll_main_shiftr1017_in[19], zll_main_shiftr1017_in[18], zll_main_shiftr1017_in[17], zll_main_shiftr1017_in[16], zll_main_shiftr1017_in[15], zll_main_shiftr1017_in[13], zll_main_shiftr1017_in[12], zll_main_shiftr1017_in[11], zll_main_shiftr1017_in[10], zll_main_shiftr1017_in[9], zll_main_shiftr1017_in[8], zll_main_shiftr1017_in[7], zll_main_shiftr1017_in[6], zll_main_shiftr1017_in[5], zll_main_shiftr1017_in[4], zll_main_shiftr1017_in[3], zll_main_shiftr1017_in[2], zll_main_shiftr1017_in[1], zll_main_shiftr1017_in[0]};
  assign zll_main_shiftr1022_in = {zll_main_shiftr1012_in[31], zll_main_shiftr1012_in[30], zll_main_shiftr1012_in[29], zll_main_shiftr1012_in[28], zll_main_shiftr1012_in[27], zll_main_shiftr1012_in[26], zll_main_shiftr1012_in[25], zll_main_shiftr1012_in[24], zll_main_shiftr1012_in[23], zll_main_shiftr1012_in[22], zll_main_shiftr1012_in[13], zll_main_shiftr1012_in[21], zll_main_shiftr1012_in[20], zll_main_shiftr1012_in[19], zll_main_shiftr1012_in[18], zll_main_shiftr1012_in[17], zll_main_shiftr1012_in[16], zll_main_shiftr1012_in[15], zll_main_shiftr1012_in[14], zll_main_shiftr1012_in[12], zll_main_shiftr1012_in[11], zll_main_shiftr1012_in[10], zll_main_shiftr1012_in[9], zll_main_shiftr1012_in[8], zll_main_shiftr1012_in[7], zll_main_shiftr1012_in[6], zll_main_shiftr1012_in[5], zll_main_shiftr1012_in[4], zll_main_shiftr1012_in[3], zll_main_shiftr1012_in[2], zll_main_shiftr1012_in[1], zll_main_shiftr1012_in[0]};
  assign zll_main_shiftr1030_in = {zll_main_shiftr1022_in[31], zll_main_shiftr1022_in[30], zll_main_shiftr1022_in[29], zll_main_shiftr1022_in[28], zll_main_shiftr1022_in[27], zll_main_shiftr1022_in[26], zll_main_shiftr1022_in[25], zll_main_shiftr1022_in[24], zll_main_shiftr1022_in[23], zll_main_shiftr1022_in[22], zll_main_shiftr1022_in[21], zll_main_shiftr1022_in[12], zll_main_shiftr1022_in[20], zll_main_shiftr1022_in[19], zll_main_shiftr1022_in[18], zll_main_shiftr1022_in[17], zll_main_shiftr1022_in[16], zll_main_shiftr1022_in[15], zll_main_shiftr1022_in[14], zll_main_shiftr1022_in[13], zll_main_shiftr1022_in[11], zll_main_shiftr1022_in[10], zll_main_shiftr1022_in[9], zll_main_shiftr1022_in[8], zll_main_shiftr1022_in[7], zll_main_shiftr1022_in[6], zll_main_shiftr1022_in[5], zll_main_shiftr1022_in[4], zll_main_shiftr1022_in[3], zll_main_shiftr1022_in[2], zll_main_shiftr1022_in[1], zll_main_shiftr1022_in[0]};
  assign zll_main_shiftr104_in = {zll_main_shiftr1030_in[31], zll_main_shiftr1030_in[30], zll_main_shiftr1030_in[29], zll_main_shiftr1030_in[11], zll_main_shiftr1030_in[28], zll_main_shiftr1030_in[27], zll_main_shiftr1030_in[26], zll_main_shiftr1030_in[25], zll_main_shiftr1030_in[24], zll_main_shiftr1030_in[23], zll_main_shiftr1030_in[22], zll_main_shiftr1030_in[21], zll_main_shiftr1030_in[20], zll_main_shiftr1030_in[19], zll_main_shiftr1030_in[18], zll_main_shiftr1030_in[17], zll_main_shiftr1030_in[16], zll_main_shiftr1030_in[15], zll_main_shiftr1030_in[14], zll_main_shiftr1030_in[13], zll_main_shiftr1030_in[12], zll_main_shiftr1030_in[10], zll_main_shiftr1030_in[9], zll_main_shiftr1030_in[8], zll_main_shiftr1030_in[7], zll_main_shiftr1030_in[6], zll_main_shiftr1030_in[5], zll_main_shiftr1030_in[4], zll_main_shiftr1030_in[3], zll_main_shiftr1030_in[2], zll_main_shiftr1030_in[1], zll_main_shiftr1030_in[0]};
  assign zll_main_shiftr1018_in = {zll_main_shiftr104_in[31], zll_main_shiftr104_in[30], zll_main_shiftr104_in[29], zll_main_shiftr104_in[28], zll_main_shiftr104_in[27], zll_main_shiftr104_in[26], zll_main_shiftr104_in[25], zll_main_shiftr104_in[10], zll_main_shiftr104_in[24], zll_main_shiftr104_in[23], zll_main_shiftr104_in[22], zll_main_shiftr104_in[21], zll_main_shiftr104_in[20], zll_main_shiftr104_in[19], zll_main_shiftr104_in[18], zll_main_shiftr104_in[17], zll_main_shiftr104_in[16], zll_main_shiftr104_in[15], zll_main_shiftr104_in[14], zll_main_shiftr104_in[13], zll_main_shiftr104_in[12], zll_main_shiftr104_in[11], zll_main_shiftr104_in[9], zll_main_shiftr104_in[8], zll_main_shiftr104_in[7], zll_main_shiftr104_in[6], zll_main_shiftr104_in[5], zll_main_shiftr104_in[4], zll_main_shiftr104_in[3], zll_main_shiftr104_in[2], zll_main_shiftr104_in[1], zll_main_shiftr104_in[0]};
  assign zll_main_shiftr1020_in = {zll_main_shiftr1018_in[31], zll_main_shiftr1018_in[30], zll_main_shiftr1018_in[29], zll_main_shiftr1018_in[28], zll_main_shiftr1018_in[27], zll_main_shiftr1018_in[26], zll_main_shiftr1018_in[25], zll_main_shiftr1018_in[24], zll_main_shiftr1018_in[23], zll_main_shiftr1018_in[22], zll_main_shiftr1018_in[21], zll_main_shiftr1018_in[20], zll_main_shiftr1018_in[19], zll_main_shiftr1018_in[18], zll_main_shiftr1018_in[17], zll_main_shiftr1018_in[16], zll_main_shiftr1018_in[15], zll_main_shiftr1018_in[14], zll_main_shiftr1018_in[13], zll_main_shiftr1018_in[12], zll_main_shiftr1018_in[11], zll_main_shiftr1018_in[10], zll_main_shiftr1018_in[8], zll_main_shiftr1018_in[7], zll_main_shiftr1018_in[6], zll_main_shiftr1018_in[5], zll_main_shiftr1018_in[4], zll_main_shiftr1018_in[3], zll_main_shiftr1018_in[2], zll_main_shiftr1018_in[1], zll_main_shiftr1018_in[0]};
  assign zll_main_shiftr107_in = {zll_main_shiftr1020_in[30], zll_main_shiftr1020_in[29], zll_main_shiftr1020_in[28], zll_main_shiftr1020_in[27], zll_main_shiftr1020_in[26], zll_main_shiftr1020_in[25], zll_main_shiftr1020_in[24], zll_main_shiftr1020_in[23], zll_main_shiftr1020_in[22], zll_main_shiftr1020_in[21], zll_main_shiftr1020_in[20], zll_main_shiftr1020_in[19], zll_main_shiftr1020_in[18], zll_main_shiftr1020_in[17], zll_main_shiftr1020_in[16], zll_main_shiftr1020_in[15], zll_main_shiftr1020_in[14], zll_main_shiftr1020_in[13], zll_main_shiftr1020_in[12], zll_main_shiftr1020_in[11], zll_main_shiftr1020_in[10], zll_main_shiftr1020_in[9], zll_main_shiftr1020_in[7], zll_main_shiftr1020_in[6], zll_main_shiftr1020_in[5], zll_main_shiftr1020_in[4], zll_main_shiftr1020_in[3], zll_main_shiftr1020_in[2], zll_main_shiftr1020_in[1], zll_main_shiftr1020_in[0]};
  assign zll_main_shiftr1027_in = {zll_main_shiftr107_in[29], zll_main_shiftr107_in[28], zll_main_shiftr107_in[27], zll_main_shiftr107_in[26], zll_main_shiftr107_in[25], zll_main_shiftr107_in[24], zll_main_shiftr107_in[23], zll_main_shiftr107_in[22], zll_main_shiftr107_in[21], zll_main_shiftr107_in[20], zll_main_shiftr107_in[19], zll_main_shiftr107_in[18], zll_main_shiftr107_in[17], zll_main_shiftr107_in[16], zll_main_shiftr107_in[15], zll_main_shiftr107_in[14], zll_main_shiftr107_in[13], zll_main_shiftr107_in[12], zll_main_shiftr107_in[11], zll_main_shiftr107_in[10], zll_main_shiftr107_in[9], zll_main_shiftr107_in[8], zll_main_shiftr107_in[6], zll_main_shiftr107_in[5], zll_main_shiftr107_in[4], zll_main_shiftr107_in[3], zll_main_shiftr107_in[2], zll_main_shiftr107_in[1], zll_main_shiftr107_in[0]};
  assign zll_main_shiftr1026_in = {zll_main_shiftr1027_in[28], zll_main_shiftr1027_in[27], zll_main_shiftr1027_in[26], zll_main_shiftr1027_in[25], zll_main_shiftr1027_in[24], zll_main_shiftr1027_in[23], zll_main_shiftr1027_in[22], zll_main_shiftr1027_in[21], zll_main_shiftr1027_in[20], zll_main_shiftr1027_in[19], zll_main_shiftr1027_in[18], zll_main_shiftr1027_in[17], zll_main_shiftr1027_in[16], zll_main_shiftr1027_in[15], zll_main_shiftr1027_in[14], zll_main_shiftr1027_in[13], zll_main_shiftr1027_in[12], zll_main_shiftr1027_in[11], zll_main_shiftr1027_in[10], zll_main_shiftr1027_in[9], zll_main_shiftr1027_in[8], zll_main_shiftr1027_in[7], zll_main_shiftr1027_in[5], zll_main_shiftr1027_in[4], zll_main_shiftr1027_in[3], zll_main_shiftr1027_in[2], zll_main_shiftr1027_in[1], zll_main_shiftr1027_in[0]};
  assign zll_main_shiftr1014_in = {zll_main_shiftr1026_in[27], zll_main_shiftr1026_in[26], zll_main_shiftr1026_in[25], zll_main_shiftr1026_in[24], zll_main_shiftr1026_in[23], zll_main_shiftr1026_in[22], zll_main_shiftr1026_in[21], zll_main_shiftr1026_in[20], zll_main_shiftr1026_in[19], zll_main_shiftr1026_in[18], zll_main_shiftr1026_in[17], zll_main_shiftr1026_in[16], zll_main_shiftr1026_in[15], zll_main_shiftr1026_in[14], zll_main_shiftr1026_in[13], zll_main_shiftr1026_in[12], zll_main_shiftr1026_in[11], zll_main_shiftr1026_in[10], zll_main_shiftr1026_in[9], zll_main_shiftr1026_in[8], zll_main_shiftr1026_in[7], zll_main_shiftr1026_in[6], zll_main_shiftr1026_in[4], zll_main_shiftr1026_in[3], zll_main_shiftr1026_in[2], zll_main_shiftr1026_in[1], zll_main_shiftr1026_in[0]};
  assign zll_main_shiftr1015_in = {zll_main_shiftr1014_in[26], zll_main_shiftr1014_in[25], zll_main_shiftr1014_in[24], zll_main_shiftr1014_in[23], zll_main_shiftr1014_in[22], zll_main_shiftr1014_in[21], zll_main_shiftr1014_in[20], zll_main_shiftr1014_in[19], zll_main_shiftr1014_in[18], zll_main_shiftr1014_in[17], zll_main_shiftr1014_in[16], zll_main_shiftr1014_in[15], zll_main_shiftr1014_in[14], zll_main_shiftr1014_in[13], zll_main_shiftr1014_in[12], zll_main_shiftr1014_in[11], zll_main_shiftr1014_in[10], zll_main_shiftr1014_in[9], zll_main_shiftr1014_in[8], zll_main_shiftr1014_in[7], zll_main_shiftr1014_in[6], zll_main_shiftr1014_in[5], zll_main_shiftr1014_in[3], zll_main_shiftr1014_in[2], zll_main_shiftr1014_in[1], zll_main_shiftr1014_in[0]};
  assign zll_main_shiftr1023_in = {zll_main_shiftr1015_in[25], zll_main_shiftr1015_in[24], zll_main_shiftr1015_in[23], zll_main_shiftr1015_in[22], zll_main_shiftr1015_in[21], zll_main_shiftr1015_in[20], zll_main_shiftr1015_in[19], zll_main_shiftr1015_in[18], zll_main_shiftr1015_in[17], zll_main_shiftr1015_in[16], zll_main_shiftr1015_in[15], zll_main_shiftr1015_in[14], zll_main_shiftr1015_in[13], zll_main_shiftr1015_in[12], zll_main_shiftr1015_in[11], zll_main_shiftr1015_in[10], zll_main_shiftr1015_in[9], zll_main_shiftr1015_in[8], zll_main_shiftr1015_in[7], zll_main_shiftr1015_in[6], zll_main_shiftr1015_in[5], zll_main_shiftr1015_in[4], zll_main_shiftr1015_in[2], zll_main_shiftr1015_in[1], zll_main_shiftr1015_in[0]};
  assign zll_main_shiftr1010_in = {zll_main_shiftr1023_in[24], zll_main_shiftr1023_in[23], zll_main_shiftr1023_in[22], zll_main_shiftr1023_in[21], zll_main_shiftr1023_in[20], zll_main_shiftr1023_in[19], zll_main_shiftr1023_in[18], zll_main_shiftr1023_in[17], zll_main_shiftr1023_in[16], zll_main_shiftr1023_in[15], zll_main_shiftr1023_in[14], zll_main_shiftr1023_in[13], zll_main_shiftr1023_in[12], zll_main_shiftr1023_in[11], zll_main_shiftr1023_in[10], zll_main_shiftr1023_in[9], zll_main_shiftr1023_in[8], zll_main_shiftr1023_in[7], zll_main_shiftr1023_in[6], zll_main_shiftr1023_in[5], zll_main_shiftr1023_in[4], zll_main_shiftr1023_in[3], zll_main_shiftr1023_in[1], zll_main_shiftr1023_in[0]};
  assign zll_main_shiftr101_in = {zll_main_shiftr1010_in[23], zll_main_shiftr1010_in[22], zll_main_shiftr1010_in[21], zll_main_shiftr1010_in[20], zll_main_shiftr1010_in[19], zll_main_shiftr1010_in[18], zll_main_shiftr1010_in[17], zll_main_shiftr1010_in[16], zll_main_shiftr1010_in[15], zll_main_shiftr1010_in[14], zll_main_shiftr1010_in[13], zll_main_shiftr1010_in[12], zll_main_shiftr1010_in[11], zll_main_shiftr1010_in[10], zll_main_shiftr1010_in[9], zll_main_shiftr1010_in[8], zll_main_shiftr1010_in[7], zll_main_shiftr1010_in[6], zll_main_shiftr1010_in[5], zll_main_shiftr1010_in[4], zll_main_shiftr1010_in[3], zll_main_shiftr1010_in[2], zll_main_shiftr1010_in[0]};
  assign xorw32_inR1 = {extres, {10'h0, zll_main_shiftr101_in[18], zll_main_shiftr101_in[14], zll_main_shiftr101_in[21], zll_main_shiftr101_in[8], zll_main_shiftr101_in[11], zll_main_shiftr101_in[20], zll_main_shiftr101_in[3], zll_main_shiftr101_in[17], zll_main_shiftr101_in[1], zll_main_shiftr101_in[5], zll_main_shiftr101_in[12], zll_main_shiftr101_in[4], zll_main_shiftr101_in[7], zll_main_shiftr101_in[22], zll_main_shiftr101_in[2], zll_main_shiftr101_in[6], zll_main_shiftr101_in[13], zll_main_shiftr101_in[16], zll_main_shiftr101_in[10], zll_main_shiftr101_in[9], zll_main_shiftr101_in[19], zll_main_shiftr101_in[15]}};
  xorW32  instR1 (xorw32_inR1[63:32], xorw32_inR1[31:0], extresR1[31:0]);
  assign plusw32_in = {extresR1, zll_main_updatesched2_in[415:384]};
  plusW32  instR2 (plusw32_in[63:32], plusw32_in[31:0], extresR2[31:0]);
  assign main_sigma0_in = zll_main_updatesched2_in[383:352];
  assign main_rotater7_in = main_sigma0_in[31:0];
  assign zll_main_rotater713_in = main_rotater7_in[31:0];
  assign zll_main_rotater7_in = {zll_main_rotater713_in[31], zll_main_rotater713_in[28], zll_main_rotater713_in[30], zll_main_rotater713_in[29], zll_main_rotater713_in[27], zll_main_rotater713_in[26], zll_main_rotater713_in[25], zll_main_rotater713_in[24], zll_main_rotater713_in[23], zll_main_rotater713_in[22], zll_main_rotater713_in[21], zll_main_rotater713_in[20], zll_main_rotater713_in[19], zll_main_rotater713_in[18], zll_main_rotater713_in[17], zll_main_rotater713_in[16], zll_main_rotater713_in[15], zll_main_rotater713_in[14], zll_main_rotater713_in[13], zll_main_rotater713_in[12], zll_main_rotater713_in[11], zll_main_rotater713_in[10], zll_main_rotater713_in[9], zll_main_rotater713_in[8], zll_main_rotater713_in[7], zll_main_rotater713_in[6], zll_main_rotater713_in[5], zll_main_rotater713_in[4], zll_main_rotater713_in[3], zll_main_rotater713_in[2], zll_main_rotater713_in[1], zll_main_rotater713_in[0]};
  assign zll_main_rotater727_in = {zll_main_rotater7_in[31], zll_main_rotater7_in[30], zll_main_rotater7_in[27], zll_main_rotater7_in[29], zll_main_rotater7_in[28], zll_main_rotater7_in[26], zll_main_rotater7_in[25], zll_main_rotater7_in[24], zll_main_rotater7_in[23], zll_main_rotater7_in[22], zll_main_rotater7_in[21], zll_main_rotater7_in[20], zll_main_rotater7_in[19], zll_main_rotater7_in[18], zll_main_rotater7_in[17], zll_main_rotater7_in[16], zll_main_rotater7_in[15], zll_main_rotater7_in[14], zll_main_rotater7_in[13], zll_main_rotater7_in[12], zll_main_rotater7_in[11], zll_main_rotater7_in[10], zll_main_rotater7_in[9], zll_main_rotater7_in[8], zll_main_rotater7_in[7], zll_main_rotater7_in[6], zll_main_rotater7_in[5], zll_main_rotater7_in[4], zll_main_rotater7_in[3], zll_main_rotater7_in[2], zll_main_rotater7_in[1], zll_main_rotater7_in[0]};
  assign zll_main_rotater76_in = {zll_main_rotater727_in[31], zll_main_rotater727_in[26], zll_main_rotater727_in[30], zll_main_rotater727_in[29], zll_main_rotater727_in[28], zll_main_rotater727_in[27], zll_main_rotater727_in[25], zll_main_rotater727_in[24], zll_main_rotater727_in[23], zll_main_rotater727_in[22], zll_main_rotater727_in[21], zll_main_rotater727_in[20], zll_main_rotater727_in[19], zll_main_rotater727_in[18], zll_main_rotater727_in[17], zll_main_rotater727_in[16], zll_main_rotater727_in[15], zll_main_rotater727_in[14], zll_main_rotater727_in[13], zll_main_rotater727_in[12], zll_main_rotater727_in[11], zll_main_rotater727_in[10], zll_main_rotater727_in[9], zll_main_rotater727_in[8], zll_main_rotater727_in[7], zll_main_rotater727_in[6], zll_main_rotater727_in[5], zll_main_rotater727_in[4], zll_main_rotater727_in[3], zll_main_rotater727_in[2], zll_main_rotater727_in[1], zll_main_rotater727_in[0]};
  assign zll_main_rotater722_in = {zll_main_rotater76_in[31], zll_main_rotater76_in[30], zll_main_rotater76_in[29], zll_main_rotater76_in[28], zll_main_rotater76_in[25], zll_main_rotater76_in[27], zll_main_rotater76_in[26], zll_main_rotater76_in[24], zll_main_rotater76_in[23], zll_main_rotater76_in[22], zll_main_rotater76_in[21], zll_main_rotater76_in[20], zll_main_rotater76_in[19], zll_main_rotater76_in[18], zll_main_rotater76_in[17], zll_main_rotater76_in[16], zll_main_rotater76_in[15], zll_main_rotater76_in[14], zll_main_rotater76_in[13], zll_main_rotater76_in[12], zll_main_rotater76_in[11], zll_main_rotater76_in[10], zll_main_rotater76_in[9], zll_main_rotater76_in[8], zll_main_rotater76_in[7], zll_main_rotater76_in[6], zll_main_rotater76_in[5], zll_main_rotater76_in[4], zll_main_rotater76_in[3], zll_main_rotater76_in[2], zll_main_rotater76_in[1], zll_main_rotater76_in[0]};
  assign zll_main_rotater725_in = {zll_main_rotater722_in[31], zll_main_rotater722_in[30], zll_main_rotater722_in[29], zll_main_rotater722_in[28], zll_main_rotater722_in[24], zll_main_rotater722_in[27], zll_main_rotater722_in[26], zll_main_rotater722_in[25], zll_main_rotater722_in[23], zll_main_rotater722_in[22], zll_main_rotater722_in[21], zll_main_rotater722_in[20], zll_main_rotater722_in[19], zll_main_rotater722_in[18], zll_main_rotater722_in[17], zll_main_rotater722_in[16], zll_main_rotater722_in[15], zll_main_rotater722_in[14], zll_main_rotater722_in[13], zll_main_rotater722_in[12], zll_main_rotater722_in[11], zll_main_rotater722_in[10], zll_main_rotater722_in[9], zll_main_rotater722_in[8], zll_main_rotater722_in[7], zll_main_rotater722_in[6], zll_main_rotater722_in[5], zll_main_rotater722_in[4], zll_main_rotater722_in[3], zll_main_rotater722_in[2], zll_main_rotater722_in[1], zll_main_rotater722_in[0]};
  assign zll_main_rotater71_in = {zll_main_rotater725_in[31], zll_main_rotater725_in[30], zll_main_rotater725_in[29], zll_main_rotater725_in[23], zll_main_rotater725_in[28], zll_main_rotater725_in[27], zll_main_rotater725_in[26], zll_main_rotater725_in[25], zll_main_rotater725_in[24], zll_main_rotater725_in[22], zll_main_rotater725_in[21], zll_main_rotater725_in[20], zll_main_rotater725_in[19], zll_main_rotater725_in[18], zll_main_rotater725_in[17], zll_main_rotater725_in[16], zll_main_rotater725_in[15], zll_main_rotater725_in[14], zll_main_rotater725_in[13], zll_main_rotater725_in[12], zll_main_rotater725_in[11], zll_main_rotater725_in[10], zll_main_rotater725_in[9], zll_main_rotater725_in[8], zll_main_rotater725_in[7], zll_main_rotater725_in[6], zll_main_rotater725_in[5], zll_main_rotater725_in[4], zll_main_rotater725_in[3], zll_main_rotater725_in[2], zll_main_rotater725_in[1], zll_main_rotater725_in[0]};
  assign zll_main_rotater75_in = {zll_main_rotater71_in[31], zll_main_rotater71_in[30], zll_main_rotater71_in[29], zll_main_rotater71_in[28], zll_main_rotater71_in[27], zll_main_rotater71_in[26], zll_main_rotater71_in[22], zll_main_rotater71_in[25], zll_main_rotater71_in[24], zll_main_rotater71_in[23], zll_main_rotater71_in[21], zll_main_rotater71_in[20], zll_main_rotater71_in[19], zll_main_rotater71_in[18], zll_main_rotater71_in[17], zll_main_rotater71_in[16], zll_main_rotater71_in[15], zll_main_rotater71_in[14], zll_main_rotater71_in[13], zll_main_rotater71_in[12], zll_main_rotater71_in[11], zll_main_rotater71_in[10], zll_main_rotater71_in[9], zll_main_rotater71_in[8], zll_main_rotater71_in[7], zll_main_rotater71_in[6], zll_main_rotater71_in[5], zll_main_rotater71_in[4], zll_main_rotater71_in[3], zll_main_rotater71_in[2], zll_main_rotater71_in[1], zll_main_rotater71_in[0]};
  assign zll_main_rotater719_in = {zll_main_rotater75_in[31], zll_main_rotater75_in[30], zll_main_rotater75_in[29], zll_main_rotater75_in[21], zll_main_rotater75_in[28], zll_main_rotater75_in[27], zll_main_rotater75_in[26], zll_main_rotater75_in[25], zll_main_rotater75_in[24], zll_main_rotater75_in[23], zll_main_rotater75_in[22], zll_main_rotater75_in[20], zll_main_rotater75_in[19], zll_main_rotater75_in[18], zll_main_rotater75_in[17], zll_main_rotater75_in[16], zll_main_rotater75_in[15], zll_main_rotater75_in[14], zll_main_rotater75_in[13], zll_main_rotater75_in[12], zll_main_rotater75_in[11], zll_main_rotater75_in[10], zll_main_rotater75_in[9], zll_main_rotater75_in[8], zll_main_rotater75_in[7], zll_main_rotater75_in[6], zll_main_rotater75_in[5], zll_main_rotater75_in[4], zll_main_rotater75_in[3], zll_main_rotater75_in[2], zll_main_rotater75_in[1], zll_main_rotater75_in[0]};
  assign zll_main_rotater728_in = {zll_main_rotater719_in[31], zll_main_rotater719_in[30], zll_main_rotater719_in[29], zll_main_rotater719_in[20], zll_main_rotater719_in[28], zll_main_rotater719_in[27], zll_main_rotater719_in[26], zll_main_rotater719_in[25], zll_main_rotater719_in[24], zll_main_rotater719_in[23], zll_main_rotater719_in[22], zll_main_rotater719_in[21], zll_main_rotater719_in[19], zll_main_rotater719_in[18], zll_main_rotater719_in[17], zll_main_rotater719_in[16], zll_main_rotater719_in[15], zll_main_rotater719_in[14], zll_main_rotater719_in[13], zll_main_rotater719_in[12], zll_main_rotater719_in[11], zll_main_rotater719_in[10], zll_main_rotater719_in[9], zll_main_rotater719_in[8], zll_main_rotater719_in[7], zll_main_rotater719_in[6], zll_main_rotater719_in[5], zll_main_rotater719_in[4], zll_main_rotater719_in[3], zll_main_rotater719_in[2], zll_main_rotater719_in[1], zll_main_rotater719_in[0]};
  assign zll_main_rotater717_in = {zll_main_rotater728_in[31], zll_main_rotater728_in[30], zll_main_rotater728_in[29], zll_main_rotater728_in[28], zll_main_rotater728_in[27], zll_main_rotater728_in[26], zll_main_rotater728_in[19], zll_main_rotater728_in[25], zll_main_rotater728_in[24], zll_main_rotater728_in[23], zll_main_rotater728_in[22], zll_main_rotater728_in[21], zll_main_rotater728_in[20], zll_main_rotater728_in[18], zll_main_rotater728_in[17], zll_main_rotater728_in[16], zll_main_rotater728_in[15], zll_main_rotater728_in[14], zll_main_rotater728_in[13], zll_main_rotater728_in[12], zll_main_rotater728_in[11], zll_main_rotater728_in[10], zll_main_rotater728_in[9], zll_main_rotater728_in[8], zll_main_rotater728_in[7], zll_main_rotater728_in[6], zll_main_rotater728_in[5], zll_main_rotater728_in[4], zll_main_rotater728_in[3], zll_main_rotater728_in[2], zll_main_rotater728_in[1], zll_main_rotater728_in[0]};
  assign zll_main_rotater731_in = {zll_main_rotater717_in[31], zll_main_rotater717_in[18], zll_main_rotater717_in[30], zll_main_rotater717_in[29], zll_main_rotater717_in[28], zll_main_rotater717_in[27], zll_main_rotater717_in[26], zll_main_rotater717_in[25], zll_main_rotater717_in[24], zll_main_rotater717_in[23], zll_main_rotater717_in[22], zll_main_rotater717_in[21], zll_main_rotater717_in[20], zll_main_rotater717_in[19], zll_main_rotater717_in[17], zll_main_rotater717_in[16], zll_main_rotater717_in[15], zll_main_rotater717_in[14], zll_main_rotater717_in[13], zll_main_rotater717_in[12], zll_main_rotater717_in[11], zll_main_rotater717_in[10], zll_main_rotater717_in[9], zll_main_rotater717_in[8], zll_main_rotater717_in[7], zll_main_rotater717_in[6], zll_main_rotater717_in[5], zll_main_rotater717_in[4], zll_main_rotater717_in[3], zll_main_rotater717_in[2], zll_main_rotater717_in[1], zll_main_rotater717_in[0]};
  assign zll_main_rotater724_in = {zll_main_rotater731_in[31], zll_main_rotater731_in[30], zll_main_rotater731_in[29], zll_main_rotater731_in[28], zll_main_rotater731_in[27], zll_main_rotater731_in[26], zll_main_rotater731_in[25], zll_main_rotater731_in[24], zll_main_rotater731_in[17], zll_main_rotater731_in[23], zll_main_rotater731_in[22], zll_main_rotater731_in[21], zll_main_rotater731_in[20], zll_main_rotater731_in[19], zll_main_rotater731_in[18], zll_main_rotater731_in[16], zll_main_rotater731_in[15], zll_main_rotater731_in[14], zll_main_rotater731_in[13], zll_main_rotater731_in[12], zll_main_rotater731_in[11], zll_main_rotater731_in[10], zll_main_rotater731_in[9], zll_main_rotater731_in[8], zll_main_rotater731_in[7], zll_main_rotater731_in[6], zll_main_rotater731_in[5], zll_main_rotater731_in[4], zll_main_rotater731_in[3], zll_main_rotater731_in[2], zll_main_rotater731_in[1], zll_main_rotater731_in[0]};
  assign zll_main_rotater711_in = {zll_main_rotater724_in[31], zll_main_rotater724_in[30], zll_main_rotater724_in[29], zll_main_rotater724_in[28], zll_main_rotater724_in[16], zll_main_rotater724_in[27], zll_main_rotater724_in[26], zll_main_rotater724_in[25], zll_main_rotater724_in[24], zll_main_rotater724_in[23], zll_main_rotater724_in[22], zll_main_rotater724_in[21], zll_main_rotater724_in[20], zll_main_rotater724_in[19], zll_main_rotater724_in[18], zll_main_rotater724_in[17], zll_main_rotater724_in[15], zll_main_rotater724_in[14], zll_main_rotater724_in[13], zll_main_rotater724_in[12], zll_main_rotater724_in[11], zll_main_rotater724_in[10], zll_main_rotater724_in[9], zll_main_rotater724_in[8], zll_main_rotater724_in[7], zll_main_rotater724_in[6], zll_main_rotater724_in[5], zll_main_rotater724_in[4], zll_main_rotater724_in[3], zll_main_rotater724_in[2], zll_main_rotater724_in[1], zll_main_rotater724_in[0]};
  assign zll_main_rotater72_in = {zll_main_rotater711_in[31], zll_main_rotater711_in[30], zll_main_rotater711_in[29], zll_main_rotater711_in[28], zll_main_rotater711_in[27], zll_main_rotater711_in[26], zll_main_rotater711_in[25], zll_main_rotater711_in[24], zll_main_rotater711_in[23], zll_main_rotater711_in[15], zll_main_rotater711_in[22], zll_main_rotater711_in[21], zll_main_rotater711_in[20], zll_main_rotater711_in[19], zll_main_rotater711_in[18], zll_main_rotater711_in[17], zll_main_rotater711_in[16], zll_main_rotater711_in[14], zll_main_rotater711_in[13], zll_main_rotater711_in[12], zll_main_rotater711_in[11], zll_main_rotater711_in[10], zll_main_rotater711_in[9], zll_main_rotater711_in[8], zll_main_rotater711_in[7], zll_main_rotater711_in[6], zll_main_rotater711_in[5], zll_main_rotater711_in[4], zll_main_rotater711_in[3], zll_main_rotater711_in[2], zll_main_rotater711_in[1], zll_main_rotater711_in[0]};
  assign zll_main_rotater720_in = {zll_main_rotater72_in[31], zll_main_rotater72_in[30], zll_main_rotater72_in[14], zll_main_rotater72_in[29], zll_main_rotater72_in[28], zll_main_rotater72_in[27], zll_main_rotater72_in[26], zll_main_rotater72_in[25], zll_main_rotater72_in[24], zll_main_rotater72_in[23], zll_main_rotater72_in[22], zll_main_rotater72_in[21], zll_main_rotater72_in[20], zll_main_rotater72_in[19], zll_main_rotater72_in[18], zll_main_rotater72_in[17], zll_main_rotater72_in[16], zll_main_rotater72_in[15], zll_main_rotater72_in[13], zll_main_rotater72_in[12], zll_main_rotater72_in[11], zll_main_rotater72_in[10], zll_main_rotater72_in[9], zll_main_rotater72_in[8], zll_main_rotater72_in[7], zll_main_rotater72_in[6], zll_main_rotater72_in[5], zll_main_rotater72_in[4], zll_main_rotater72_in[3], zll_main_rotater72_in[2], zll_main_rotater72_in[1], zll_main_rotater72_in[0]};
  assign zll_main_rotater718_in = {zll_main_rotater720_in[31], zll_main_rotater720_in[30], zll_main_rotater720_in[29], zll_main_rotater720_in[28], zll_main_rotater720_in[27], zll_main_rotater720_in[26], zll_main_rotater720_in[25], zll_main_rotater720_in[24], zll_main_rotater720_in[23], zll_main_rotater720_in[22], zll_main_rotater720_in[21], zll_main_rotater720_in[20], zll_main_rotater720_in[19], zll_main_rotater720_in[18], zll_main_rotater720_in[17], zll_main_rotater720_in[16], zll_main_rotater720_in[15], zll_main_rotater720_in[13], zll_main_rotater720_in[14], zll_main_rotater720_in[12], zll_main_rotater720_in[11], zll_main_rotater720_in[10], zll_main_rotater720_in[9], zll_main_rotater720_in[8], zll_main_rotater720_in[7], zll_main_rotater720_in[6], zll_main_rotater720_in[5], zll_main_rotater720_in[4], zll_main_rotater720_in[3], zll_main_rotater720_in[2], zll_main_rotater720_in[1], zll_main_rotater720_in[0]};
  assign zll_main_rotater79_in = {zll_main_rotater718_in[31], zll_main_rotater718_in[30], zll_main_rotater718_in[29], zll_main_rotater718_in[28], zll_main_rotater718_in[27], zll_main_rotater718_in[26], zll_main_rotater718_in[25], zll_main_rotater718_in[24], zll_main_rotater718_in[23], zll_main_rotater718_in[22], zll_main_rotater718_in[21], zll_main_rotater718_in[20], zll_main_rotater718_in[19], zll_main_rotater718_in[18], zll_main_rotater718_in[17], zll_main_rotater718_in[16], zll_main_rotater718_in[15], zll_main_rotater718_in[12], zll_main_rotater718_in[14], zll_main_rotater718_in[13], zll_main_rotater718_in[11], zll_main_rotater718_in[10], zll_main_rotater718_in[9], zll_main_rotater718_in[8], zll_main_rotater718_in[7], zll_main_rotater718_in[6], zll_main_rotater718_in[5], zll_main_rotater718_in[4], zll_main_rotater718_in[3], zll_main_rotater718_in[2], zll_main_rotater718_in[1], zll_main_rotater718_in[0]};
  assign zll_main_rotater714_in = {zll_main_rotater79_in[31], zll_main_rotater79_in[30], zll_main_rotater79_in[29], zll_main_rotater79_in[28], zll_main_rotater79_in[27], zll_main_rotater79_in[26], zll_main_rotater79_in[25], zll_main_rotater79_in[24], zll_main_rotater79_in[23], zll_main_rotater79_in[22], zll_main_rotater79_in[21], zll_main_rotater79_in[20], zll_main_rotater79_in[11], zll_main_rotater79_in[19], zll_main_rotater79_in[18], zll_main_rotater79_in[17], zll_main_rotater79_in[16], zll_main_rotater79_in[15], zll_main_rotater79_in[14], zll_main_rotater79_in[13], zll_main_rotater79_in[12], zll_main_rotater79_in[10], zll_main_rotater79_in[9], zll_main_rotater79_in[8], zll_main_rotater79_in[7], zll_main_rotater79_in[6], zll_main_rotater79_in[5], zll_main_rotater79_in[4], zll_main_rotater79_in[3], zll_main_rotater79_in[2], zll_main_rotater79_in[1], zll_main_rotater79_in[0]};
  assign zll_main_rotater74_in = {zll_main_rotater714_in[31], zll_main_rotater714_in[30], zll_main_rotater714_in[29], zll_main_rotater714_in[28], zll_main_rotater714_in[27], zll_main_rotater714_in[26], zll_main_rotater714_in[25], zll_main_rotater714_in[24], zll_main_rotater714_in[23], zll_main_rotater714_in[22], zll_main_rotater714_in[21], zll_main_rotater714_in[20], zll_main_rotater714_in[19], zll_main_rotater714_in[18], zll_main_rotater714_in[17], zll_main_rotater714_in[16], zll_main_rotater714_in[15], zll_main_rotater714_in[14], zll_main_rotater714_in[10], zll_main_rotater714_in[13], zll_main_rotater714_in[12], zll_main_rotater714_in[11], zll_main_rotater714_in[9], zll_main_rotater714_in[8], zll_main_rotater714_in[7], zll_main_rotater714_in[6], zll_main_rotater714_in[5], zll_main_rotater714_in[4], zll_main_rotater714_in[3], zll_main_rotater714_in[2], zll_main_rotater714_in[1], zll_main_rotater714_in[0]};
  assign zll_main_rotater77_in = {zll_main_rotater74_in[31], zll_main_rotater74_in[30], zll_main_rotater74_in[29], zll_main_rotater74_in[28], zll_main_rotater74_in[27], zll_main_rotater74_in[26], zll_main_rotater74_in[25], zll_main_rotater74_in[24], zll_main_rotater74_in[9], zll_main_rotater74_in[23], zll_main_rotater74_in[22], zll_main_rotater74_in[21], zll_main_rotater74_in[20], zll_main_rotater74_in[19], zll_main_rotater74_in[18], zll_main_rotater74_in[17], zll_main_rotater74_in[16], zll_main_rotater74_in[15], zll_main_rotater74_in[14], zll_main_rotater74_in[13], zll_main_rotater74_in[12], zll_main_rotater74_in[11], zll_main_rotater74_in[10], zll_main_rotater74_in[8], zll_main_rotater74_in[7], zll_main_rotater74_in[6], zll_main_rotater74_in[5], zll_main_rotater74_in[4], zll_main_rotater74_in[3], zll_main_rotater74_in[2], zll_main_rotater74_in[1], zll_main_rotater74_in[0]};
  assign zll_main_rotater712_in = {zll_main_rotater77_in[31], zll_main_rotater77_in[30], zll_main_rotater77_in[29], zll_main_rotater77_in[28], zll_main_rotater77_in[27], zll_main_rotater77_in[26], zll_main_rotater77_in[25], zll_main_rotater77_in[24], zll_main_rotater77_in[23], zll_main_rotater77_in[22], zll_main_rotater77_in[21], zll_main_rotater77_in[8], zll_main_rotater77_in[20], zll_main_rotater77_in[19], zll_main_rotater77_in[18], zll_main_rotater77_in[17], zll_main_rotater77_in[16], zll_main_rotater77_in[15], zll_main_rotater77_in[14], zll_main_rotater77_in[13], zll_main_rotater77_in[12], zll_main_rotater77_in[11], zll_main_rotater77_in[10], zll_main_rotater77_in[9], zll_main_rotater77_in[7], zll_main_rotater77_in[6], zll_main_rotater77_in[5], zll_main_rotater77_in[4], zll_main_rotater77_in[3], zll_main_rotater77_in[2], zll_main_rotater77_in[1], zll_main_rotater77_in[0]};
  assign zll_main_rotater721_in = {zll_main_rotater712_in[31], zll_main_rotater712_in[30], zll_main_rotater712_in[29], zll_main_rotater712_in[28], zll_main_rotater712_in[27], zll_main_rotater712_in[26], zll_main_rotater712_in[25], zll_main_rotater712_in[24], zll_main_rotater712_in[23], zll_main_rotater712_in[22], zll_main_rotater712_in[21], zll_main_rotater712_in[20], zll_main_rotater712_in[19], zll_main_rotater712_in[18], zll_main_rotater712_in[17], zll_main_rotater712_in[16], zll_main_rotater712_in[7], zll_main_rotater712_in[15], zll_main_rotater712_in[14], zll_main_rotater712_in[13], zll_main_rotater712_in[12], zll_main_rotater712_in[11], zll_main_rotater712_in[10], zll_main_rotater712_in[9], zll_main_rotater712_in[8], zll_main_rotater712_in[6], zll_main_rotater712_in[5], zll_main_rotater712_in[4], zll_main_rotater712_in[3], zll_main_rotater712_in[2], zll_main_rotater712_in[1], zll_main_rotater712_in[0]};
  assign zll_main_rotater729_in = {zll_main_rotater721_in[31], zll_main_rotater721_in[30], zll_main_rotater721_in[29], zll_main_rotater721_in[28], zll_main_rotater721_in[27], zll_main_rotater721_in[26], zll_main_rotater721_in[25], zll_main_rotater721_in[24], zll_main_rotater721_in[23], zll_main_rotater721_in[22], zll_main_rotater721_in[21], zll_main_rotater721_in[20], zll_main_rotater721_in[19], zll_main_rotater721_in[18], zll_main_rotater721_in[17], zll_main_rotater721_in[16], zll_main_rotater721_in[15], zll_main_rotater721_in[6], zll_main_rotater721_in[14], zll_main_rotater721_in[13], zll_main_rotater721_in[12], zll_main_rotater721_in[11], zll_main_rotater721_in[10], zll_main_rotater721_in[9], zll_main_rotater721_in[8], zll_main_rotater721_in[7], zll_main_rotater721_in[5], zll_main_rotater721_in[4], zll_main_rotater721_in[3], zll_main_rotater721_in[2], zll_main_rotater721_in[1], zll_main_rotater721_in[0]};
  assign zll_main_rotater726_in = {zll_main_rotater729_in[31], zll_main_rotater729_in[30], zll_main_rotater729_in[29], zll_main_rotater729_in[28], zll_main_rotater729_in[27], zll_main_rotater729_in[5], zll_main_rotater729_in[26], zll_main_rotater729_in[25], zll_main_rotater729_in[24], zll_main_rotater729_in[23], zll_main_rotater729_in[22], zll_main_rotater729_in[21], zll_main_rotater729_in[20], zll_main_rotater729_in[19], zll_main_rotater729_in[18], zll_main_rotater729_in[17], zll_main_rotater729_in[16], zll_main_rotater729_in[15], zll_main_rotater729_in[14], zll_main_rotater729_in[13], zll_main_rotater729_in[12], zll_main_rotater729_in[11], zll_main_rotater729_in[10], zll_main_rotater729_in[9], zll_main_rotater729_in[8], zll_main_rotater729_in[7], zll_main_rotater729_in[6], zll_main_rotater729_in[4], zll_main_rotater729_in[3], zll_main_rotater729_in[2], zll_main_rotater729_in[1], zll_main_rotater729_in[0]};
  assign zll_main_rotater73_in = {zll_main_rotater726_in[31], zll_main_rotater726_in[30], zll_main_rotater726_in[29], zll_main_rotater726_in[28], zll_main_rotater726_in[27], zll_main_rotater726_in[26], zll_main_rotater726_in[25], zll_main_rotater726_in[24], zll_main_rotater726_in[23], zll_main_rotater726_in[22], zll_main_rotater726_in[21], zll_main_rotater726_in[20], zll_main_rotater726_in[19], zll_main_rotater726_in[18], zll_main_rotater726_in[17], zll_main_rotater726_in[16], zll_main_rotater726_in[15], zll_main_rotater726_in[4], zll_main_rotater726_in[14], zll_main_rotater726_in[13], zll_main_rotater726_in[12], zll_main_rotater726_in[11], zll_main_rotater726_in[10], zll_main_rotater726_in[9], zll_main_rotater726_in[8], zll_main_rotater726_in[7], zll_main_rotater726_in[6], zll_main_rotater726_in[5], zll_main_rotater726_in[3], zll_main_rotater726_in[2], zll_main_rotater726_in[1], zll_main_rotater726_in[0]};
  assign zll_main_rotater78_in = {zll_main_rotater73_in[31], zll_main_rotater73_in[30], zll_main_rotater73_in[29], zll_main_rotater73_in[28], zll_main_rotater73_in[27], zll_main_rotater73_in[3], zll_main_rotater73_in[26], zll_main_rotater73_in[25], zll_main_rotater73_in[24], zll_main_rotater73_in[23], zll_main_rotater73_in[22], zll_main_rotater73_in[21], zll_main_rotater73_in[20], zll_main_rotater73_in[19], zll_main_rotater73_in[18], zll_main_rotater73_in[17], zll_main_rotater73_in[16], zll_main_rotater73_in[15], zll_main_rotater73_in[14], zll_main_rotater73_in[13], zll_main_rotater73_in[12], zll_main_rotater73_in[11], zll_main_rotater73_in[10], zll_main_rotater73_in[9], zll_main_rotater73_in[8], zll_main_rotater73_in[7], zll_main_rotater73_in[6], zll_main_rotater73_in[5], zll_main_rotater73_in[4], zll_main_rotater73_in[2], zll_main_rotater73_in[1], zll_main_rotater73_in[0]};
  assign zll_main_rotater716_in = {zll_main_rotater78_in[31], zll_main_rotater78_in[30], zll_main_rotater78_in[29], zll_main_rotater78_in[28], zll_main_rotater78_in[27], zll_main_rotater78_in[26], zll_main_rotater78_in[25], zll_main_rotater78_in[24], zll_main_rotater78_in[23], zll_main_rotater78_in[22], zll_main_rotater78_in[21], zll_main_rotater78_in[20], zll_main_rotater78_in[19], zll_main_rotater78_in[18], zll_main_rotater78_in[17], zll_main_rotater78_in[16], zll_main_rotater78_in[15], zll_main_rotater78_in[14], zll_main_rotater78_in[13], zll_main_rotater78_in[12], zll_main_rotater78_in[11], zll_main_rotater78_in[10], zll_main_rotater78_in[9], zll_main_rotater78_in[8], zll_main_rotater78_in[7], zll_main_rotater78_in[6], zll_main_rotater78_in[5], zll_main_rotater78_in[4], zll_main_rotater78_in[2], zll_main_rotater78_in[3], zll_main_rotater78_in[1], zll_main_rotater78_in[0]};
  assign zll_main_rotater715_in = {zll_main_rotater716_in[31], zll_main_rotater716_in[30], zll_main_rotater716_in[29], zll_main_rotater716_in[28], zll_main_rotater716_in[27], zll_main_rotater716_in[26], zll_main_rotater716_in[25], zll_main_rotater716_in[24], zll_main_rotater716_in[1], zll_main_rotater716_in[23], zll_main_rotater716_in[22], zll_main_rotater716_in[21], zll_main_rotater716_in[20], zll_main_rotater716_in[19], zll_main_rotater716_in[18], zll_main_rotater716_in[17], zll_main_rotater716_in[16], zll_main_rotater716_in[15], zll_main_rotater716_in[14], zll_main_rotater716_in[13], zll_main_rotater716_in[12], zll_main_rotater716_in[11], zll_main_rotater716_in[10], zll_main_rotater716_in[9], zll_main_rotater716_in[8], zll_main_rotater716_in[7], zll_main_rotater716_in[6], zll_main_rotater716_in[5], zll_main_rotater716_in[4], zll_main_rotater716_in[3], zll_main_rotater716_in[2], zll_main_rotater716_in[0]};
  assign main_rotater18_in = main_sigma0_in[31:0];
  assign zll_main_rotater1825_in = main_rotater18_in[31:0];
  assign zll_main_rotater1818_in = {zll_main_rotater1825_in[30], zll_main_rotater1825_in[31], zll_main_rotater1825_in[29], zll_main_rotater1825_in[28], zll_main_rotater1825_in[27], zll_main_rotater1825_in[26], zll_main_rotater1825_in[25], zll_main_rotater1825_in[24], zll_main_rotater1825_in[23], zll_main_rotater1825_in[22], zll_main_rotater1825_in[21], zll_main_rotater1825_in[20], zll_main_rotater1825_in[19], zll_main_rotater1825_in[18], zll_main_rotater1825_in[17], zll_main_rotater1825_in[16], zll_main_rotater1825_in[15], zll_main_rotater1825_in[14], zll_main_rotater1825_in[13], zll_main_rotater1825_in[12], zll_main_rotater1825_in[11], zll_main_rotater1825_in[10], zll_main_rotater1825_in[9], zll_main_rotater1825_in[8], zll_main_rotater1825_in[7], zll_main_rotater1825_in[6], zll_main_rotater1825_in[5], zll_main_rotater1825_in[4], zll_main_rotater1825_in[3], zll_main_rotater1825_in[2], zll_main_rotater1825_in[1], zll_main_rotater1825_in[0]};
  assign zll_main_rotater1828_in = {zll_main_rotater1818_in[29], zll_main_rotater1818_in[31], zll_main_rotater1818_in[30], zll_main_rotater1818_in[28], zll_main_rotater1818_in[27], zll_main_rotater1818_in[26], zll_main_rotater1818_in[25], zll_main_rotater1818_in[24], zll_main_rotater1818_in[23], zll_main_rotater1818_in[22], zll_main_rotater1818_in[21], zll_main_rotater1818_in[20], zll_main_rotater1818_in[19], zll_main_rotater1818_in[18], zll_main_rotater1818_in[17], zll_main_rotater1818_in[16], zll_main_rotater1818_in[15], zll_main_rotater1818_in[14], zll_main_rotater1818_in[13], zll_main_rotater1818_in[12], zll_main_rotater1818_in[11], zll_main_rotater1818_in[10], zll_main_rotater1818_in[9], zll_main_rotater1818_in[8], zll_main_rotater1818_in[7], zll_main_rotater1818_in[6], zll_main_rotater1818_in[5], zll_main_rotater1818_in[4], zll_main_rotater1818_in[3], zll_main_rotater1818_in[2], zll_main_rotater1818_in[1], zll_main_rotater1818_in[0]};
  assign zll_main_rotater1826_in = {zll_main_rotater1828_in[31], zll_main_rotater1828_in[30], zll_main_rotater1828_in[28], zll_main_rotater1828_in[29], zll_main_rotater1828_in[27], zll_main_rotater1828_in[26], zll_main_rotater1828_in[25], zll_main_rotater1828_in[24], zll_main_rotater1828_in[23], zll_main_rotater1828_in[22], zll_main_rotater1828_in[21], zll_main_rotater1828_in[20], zll_main_rotater1828_in[19], zll_main_rotater1828_in[18], zll_main_rotater1828_in[17], zll_main_rotater1828_in[16], zll_main_rotater1828_in[15], zll_main_rotater1828_in[14], zll_main_rotater1828_in[13], zll_main_rotater1828_in[12], zll_main_rotater1828_in[11], zll_main_rotater1828_in[10], zll_main_rotater1828_in[9], zll_main_rotater1828_in[8], zll_main_rotater1828_in[7], zll_main_rotater1828_in[6], zll_main_rotater1828_in[5], zll_main_rotater1828_in[4], zll_main_rotater1828_in[3], zll_main_rotater1828_in[2], zll_main_rotater1828_in[1], zll_main_rotater1828_in[0]};
  assign zll_main_rotater1824_in = {zll_main_rotater1826_in[27], zll_main_rotater1826_in[31], zll_main_rotater1826_in[30], zll_main_rotater1826_in[29], zll_main_rotater1826_in[28], zll_main_rotater1826_in[26], zll_main_rotater1826_in[25], zll_main_rotater1826_in[24], zll_main_rotater1826_in[23], zll_main_rotater1826_in[22], zll_main_rotater1826_in[21], zll_main_rotater1826_in[20], zll_main_rotater1826_in[19], zll_main_rotater1826_in[18], zll_main_rotater1826_in[17], zll_main_rotater1826_in[16], zll_main_rotater1826_in[15], zll_main_rotater1826_in[14], zll_main_rotater1826_in[13], zll_main_rotater1826_in[12], zll_main_rotater1826_in[11], zll_main_rotater1826_in[10], zll_main_rotater1826_in[9], zll_main_rotater1826_in[8], zll_main_rotater1826_in[7], zll_main_rotater1826_in[6], zll_main_rotater1826_in[5], zll_main_rotater1826_in[4], zll_main_rotater1826_in[3], zll_main_rotater1826_in[2], zll_main_rotater1826_in[1], zll_main_rotater1826_in[0]};
  assign zll_main_rotater188_in = {zll_main_rotater1824_in[26], zll_main_rotater1824_in[31], zll_main_rotater1824_in[30], zll_main_rotater1824_in[29], zll_main_rotater1824_in[28], zll_main_rotater1824_in[27], zll_main_rotater1824_in[25], zll_main_rotater1824_in[24], zll_main_rotater1824_in[23], zll_main_rotater1824_in[22], zll_main_rotater1824_in[21], zll_main_rotater1824_in[20], zll_main_rotater1824_in[19], zll_main_rotater1824_in[18], zll_main_rotater1824_in[17], zll_main_rotater1824_in[16], zll_main_rotater1824_in[15], zll_main_rotater1824_in[14], zll_main_rotater1824_in[13], zll_main_rotater1824_in[12], zll_main_rotater1824_in[11], zll_main_rotater1824_in[10], zll_main_rotater1824_in[9], zll_main_rotater1824_in[8], zll_main_rotater1824_in[7], zll_main_rotater1824_in[6], zll_main_rotater1824_in[5], zll_main_rotater1824_in[4], zll_main_rotater1824_in[3], zll_main_rotater1824_in[2], zll_main_rotater1824_in[1], zll_main_rotater1824_in[0]};
  assign zll_main_rotater1817_in = {zll_main_rotater188_in[31], zll_main_rotater188_in[24], zll_main_rotater188_in[30], zll_main_rotater188_in[29], zll_main_rotater188_in[28], zll_main_rotater188_in[27], zll_main_rotater188_in[26], zll_main_rotater188_in[25], zll_main_rotater188_in[23], zll_main_rotater188_in[22], zll_main_rotater188_in[21], zll_main_rotater188_in[20], zll_main_rotater188_in[19], zll_main_rotater188_in[18], zll_main_rotater188_in[17], zll_main_rotater188_in[16], zll_main_rotater188_in[15], zll_main_rotater188_in[14], zll_main_rotater188_in[13], zll_main_rotater188_in[12], zll_main_rotater188_in[11], zll_main_rotater188_in[10], zll_main_rotater188_in[9], zll_main_rotater188_in[8], zll_main_rotater188_in[7], zll_main_rotater188_in[6], zll_main_rotater188_in[5], zll_main_rotater188_in[4], zll_main_rotater188_in[3], zll_main_rotater188_in[2], zll_main_rotater188_in[1], zll_main_rotater188_in[0]};
  assign zll_main_rotater181_in = {zll_main_rotater1817_in[31], zll_main_rotater1817_in[30], zll_main_rotater1817_in[29], zll_main_rotater1817_in[28], zll_main_rotater1817_in[27], zll_main_rotater1817_in[26], zll_main_rotater1817_in[23], zll_main_rotater1817_in[25], zll_main_rotater1817_in[24], zll_main_rotater1817_in[22], zll_main_rotater1817_in[21], zll_main_rotater1817_in[20], zll_main_rotater1817_in[19], zll_main_rotater1817_in[18], zll_main_rotater1817_in[17], zll_main_rotater1817_in[16], zll_main_rotater1817_in[15], zll_main_rotater1817_in[14], zll_main_rotater1817_in[13], zll_main_rotater1817_in[12], zll_main_rotater1817_in[11], zll_main_rotater1817_in[10], zll_main_rotater1817_in[9], zll_main_rotater1817_in[8], zll_main_rotater1817_in[7], zll_main_rotater1817_in[6], zll_main_rotater1817_in[5], zll_main_rotater1817_in[4], zll_main_rotater1817_in[3], zll_main_rotater1817_in[2], zll_main_rotater1817_in[1], zll_main_rotater1817_in[0]};
  assign zll_main_rotater1811_in = {zll_main_rotater181_in[31], zll_main_rotater181_in[22], zll_main_rotater181_in[30], zll_main_rotater181_in[29], zll_main_rotater181_in[28], zll_main_rotater181_in[27], zll_main_rotater181_in[26], zll_main_rotater181_in[25], zll_main_rotater181_in[24], zll_main_rotater181_in[23], zll_main_rotater181_in[21], zll_main_rotater181_in[20], zll_main_rotater181_in[19], zll_main_rotater181_in[18], zll_main_rotater181_in[17], zll_main_rotater181_in[16], zll_main_rotater181_in[15], zll_main_rotater181_in[14], zll_main_rotater181_in[13], zll_main_rotater181_in[12], zll_main_rotater181_in[11], zll_main_rotater181_in[10], zll_main_rotater181_in[9], zll_main_rotater181_in[8], zll_main_rotater181_in[7], zll_main_rotater181_in[6], zll_main_rotater181_in[5], zll_main_rotater181_in[4], zll_main_rotater181_in[3], zll_main_rotater181_in[2], zll_main_rotater181_in[1], zll_main_rotater181_in[0]};
  assign zll_main_rotater1830_in = {zll_main_rotater1811_in[21], zll_main_rotater1811_in[31], zll_main_rotater1811_in[30], zll_main_rotater1811_in[29], zll_main_rotater1811_in[28], zll_main_rotater1811_in[27], zll_main_rotater1811_in[26], zll_main_rotater1811_in[25], zll_main_rotater1811_in[24], zll_main_rotater1811_in[23], zll_main_rotater1811_in[22], zll_main_rotater1811_in[20], zll_main_rotater1811_in[19], zll_main_rotater1811_in[18], zll_main_rotater1811_in[17], zll_main_rotater1811_in[16], zll_main_rotater1811_in[15], zll_main_rotater1811_in[14], zll_main_rotater1811_in[13], zll_main_rotater1811_in[12], zll_main_rotater1811_in[11], zll_main_rotater1811_in[10], zll_main_rotater1811_in[9], zll_main_rotater1811_in[8], zll_main_rotater1811_in[7], zll_main_rotater1811_in[6], zll_main_rotater1811_in[5], zll_main_rotater1811_in[4], zll_main_rotater1811_in[3], zll_main_rotater1811_in[2], zll_main_rotater1811_in[1], zll_main_rotater1811_in[0]};
  assign zll_main_rotater1821_in = {zll_main_rotater1830_in[31], zll_main_rotater1830_in[30], zll_main_rotater1830_in[29], zll_main_rotater1830_in[28], zll_main_rotater1830_in[27], zll_main_rotater1830_in[26], zll_main_rotater1830_in[25], zll_main_rotater1830_in[24], zll_main_rotater1830_in[23], zll_main_rotater1830_in[20], zll_main_rotater1830_in[22], zll_main_rotater1830_in[21], zll_main_rotater1830_in[19], zll_main_rotater1830_in[18], zll_main_rotater1830_in[17], zll_main_rotater1830_in[16], zll_main_rotater1830_in[15], zll_main_rotater1830_in[14], zll_main_rotater1830_in[13], zll_main_rotater1830_in[12], zll_main_rotater1830_in[11], zll_main_rotater1830_in[10], zll_main_rotater1830_in[9], zll_main_rotater1830_in[8], zll_main_rotater1830_in[7], zll_main_rotater1830_in[6], zll_main_rotater1830_in[5], zll_main_rotater1830_in[4], zll_main_rotater1830_in[3], zll_main_rotater1830_in[2], zll_main_rotater1830_in[1], zll_main_rotater1830_in[0]};
  assign zll_main_rotater1813_in = {zll_main_rotater1821_in[31], zll_main_rotater1821_in[30], zll_main_rotater1821_in[29], zll_main_rotater1821_in[28], zll_main_rotater1821_in[27], zll_main_rotater1821_in[26], zll_main_rotater1821_in[25], zll_main_rotater1821_in[19], zll_main_rotater1821_in[24], zll_main_rotater1821_in[23], zll_main_rotater1821_in[22], zll_main_rotater1821_in[21], zll_main_rotater1821_in[20], zll_main_rotater1821_in[18], zll_main_rotater1821_in[17], zll_main_rotater1821_in[16], zll_main_rotater1821_in[15], zll_main_rotater1821_in[14], zll_main_rotater1821_in[13], zll_main_rotater1821_in[12], zll_main_rotater1821_in[11], zll_main_rotater1821_in[10], zll_main_rotater1821_in[9], zll_main_rotater1821_in[8], zll_main_rotater1821_in[7], zll_main_rotater1821_in[6], zll_main_rotater1821_in[5], zll_main_rotater1821_in[4], zll_main_rotater1821_in[3], zll_main_rotater1821_in[2], zll_main_rotater1821_in[1], zll_main_rotater1821_in[0]};
  assign zll_main_rotater186_in = {zll_main_rotater1813_in[31], zll_main_rotater1813_in[30], zll_main_rotater1813_in[29], zll_main_rotater1813_in[28], zll_main_rotater1813_in[27], zll_main_rotater1813_in[26], zll_main_rotater1813_in[25], zll_main_rotater1813_in[24], zll_main_rotater1813_in[23], zll_main_rotater1813_in[22], zll_main_rotater1813_in[18], zll_main_rotater1813_in[21], zll_main_rotater1813_in[20], zll_main_rotater1813_in[19], zll_main_rotater1813_in[17], zll_main_rotater1813_in[16], zll_main_rotater1813_in[15], zll_main_rotater1813_in[14], zll_main_rotater1813_in[13], zll_main_rotater1813_in[12], zll_main_rotater1813_in[11], zll_main_rotater1813_in[10], zll_main_rotater1813_in[9], zll_main_rotater1813_in[8], zll_main_rotater1813_in[7], zll_main_rotater1813_in[6], zll_main_rotater1813_in[5], zll_main_rotater1813_in[4], zll_main_rotater1813_in[3], zll_main_rotater1813_in[2], zll_main_rotater1813_in[1], zll_main_rotater1813_in[0]};
  assign zll_main_rotater1827_in = {zll_main_rotater186_in[31], zll_main_rotater186_in[30], zll_main_rotater186_in[29], zll_main_rotater186_in[28], zll_main_rotater186_in[27], zll_main_rotater186_in[17], zll_main_rotater186_in[26], zll_main_rotater186_in[25], zll_main_rotater186_in[24], zll_main_rotater186_in[23], zll_main_rotater186_in[22], zll_main_rotater186_in[21], zll_main_rotater186_in[20], zll_main_rotater186_in[19], zll_main_rotater186_in[18], zll_main_rotater186_in[16], zll_main_rotater186_in[15], zll_main_rotater186_in[14], zll_main_rotater186_in[13], zll_main_rotater186_in[12], zll_main_rotater186_in[11], zll_main_rotater186_in[10], zll_main_rotater186_in[9], zll_main_rotater186_in[8], zll_main_rotater186_in[7], zll_main_rotater186_in[6], zll_main_rotater186_in[5], zll_main_rotater186_in[4], zll_main_rotater186_in[3], zll_main_rotater186_in[2], zll_main_rotater186_in[1], zll_main_rotater186_in[0]};
  assign zll_main_rotater185_in = {zll_main_rotater1827_in[31], zll_main_rotater1827_in[30], zll_main_rotater1827_in[16], zll_main_rotater1827_in[29], zll_main_rotater1827_in[28], zll_main_rotater1827_in[27], zll_main_rotater1827_in[26], zll_main_rotater1827_in[25], zll_main_rotater1827_in[24], zll_main_rotater1827_in[23], zll_main_rotater1827_in[22], zll_main_rotater1827_in[21], zll_main_rotater1827_in[20], zll_main_rotater1827_in[19], zll_main_rotater1827_in[18], zll_main_rotater1827_in[17], zll_main_rotater1827_in[15], zll_main_rotater1827_in[14], zll_main_rotater1827_in[13], zll_main_rotater1827_in[12], zll_main_rotater1827_in[11], zll_main_rotater1827_in[10], zll_main_rotater1827_in[9], zll_main_rotater1827_in[8], zll_main_rotater1827_in[7], zll_main_rotater1827_in[6], zll_main_rotater1827_in[5], zll_main_rotater1827_in[4], zll_main_rotater1827_in[3], zll_main_rotater1827_in[2], zll_main_rotater1827_in[1], zll_main_rotater1827_in[0]};
  assign zll_main_rotater1820_in = {zll_main_rotater185_in[31], zll_main_rotater185_in[30], zll_main_rotater185_in[29], zll_main_rotater185_in[28], zll_main_rotater185_in[27], zll_main_rotater185_in[26], zll_main_rotater185_in[25], zll_main_rotater185_in[24], zll_main_rotater185_in[23], zll_main_rotater185_in[22], zll_main_rotater185_in[21], zll_main_rotater185_in[20], zll_main_rotater185_in[15], zll_main_rotater185_in[19], zll_main_rotater185_in[18], zll_main_rotater185_in[17], zll_main_rotater185_in[16], zll_main_rotater185_in[14], zll_main_rotater185_in[13], zll_main_rotater185_in[12], zll_main_rotater185_in[11], zll_main_rotater185_in[10], zll_main_rotater185_in[9], zll_main_rotater185_in[8], zll_main_rotater185_in[7], zll_main_rotater185_in[6], zll_main_rotater185_in[5], zll_main_rotater185_in[4], zll_main_rotater185_in[3], zll_main_rotater185_in[2], zll_main_rotater185_in[1], zll_main_rotater185_in[0]};
  assign zll_main_rotater1822_in = {zll_main_rotater1820_in[31], zll_main_rotater1820_in[30], zll_main_rotater1820_in[29], zll_main_rotater1820_in[14], zll_main_rotater1820_in[28], zll_main_rotater1820_in[27], zll_main_rotater1820_in[26], zll_main_rotater1820_in[25], zll_main_rotater1820_in[24], zll_main_rotater1820_in[23], zll_main_rotater1820_in[22], zll_main_rotater1820_in[21], zll_main_rotater1820_in[20], zll_main_rotater1820_in[19], zll_main_rotater1820_in[18], zll_main_rotater1820_in[17], zll_main_rotater1820_in[16], zll_main_rotater1820_in[15], zll_main_rotater1820_in[13], zll_main_rotater1820_in[12], zll_main_rotater1820_in[11], zll_main_rotater1820_in[10], zll_main_rotater1820_in[9], zll_main_rotater1820_in[8], zll_main_rotater1820_in[7], zll_main_rotater1820_in[6], zll_main_rotater1820_in[5], zll_main_rotater1820_in[4], zll_main_rotater1820_in[3], zll_main_rotater1820_in[2], zll_main_rotater1820_in[1], zll_main_rotater1820_in[0]};
  assign zll_main_rotater1814_in = {zll_main_rotater1822_in[31], zll_main_rotater1822_in[30], zll_main_rotater1822_in[29], zll_main_rotater1822_in[28], zll_main_rotater1822_in[27], zll_main_rotater1822_in[26], zll_main_rotater1822_in[25], zll_main_rotater1822_in[24], zll_main_rotater1822_in[23], zll_main_rotater1822_in[22], zll_main_rotater1822_in[21], zll_main_rotater1822_in[20], zll_main_rotater1822_in[19], zll_main_rotater1822_in[18], zll_main_rotater1822_in[13], zll_main_rotater1822_in[17], zll_main_rotater1822_in[16], zll_main_rotater1822_in[15], zll_main_rotater1822_in[14], zll_main_rotater1822_in[12], zll_main_rotater1822_in[11], zll_main_rotater1822_in[10], zll_main_rotater1822_in[9], zll_main_rotater1822_in[8], zll_main_rotater1822_in[7], zll_main_rotater1822_in[6], zll_main_rotater1822_in[5], zll_main_rotater1822_in[4], zll_main_rotater1822_in[3], zll_main_rotater1822_in[2], zll_main_rotater1822_in[1], zll_main_rotater1822_in[0]};
  assign zll_main_rotater1815_in = {zll_main_rotater1814_in[31], zll_main_rotater1814_in[30], zll_main_rotater1814_in[29], zll_main_rotater1814_in[28], zll_main_rotater1814_in[27], zll_main_rotater1814_in[26], zll_main_rotater1814_in[25], zll_main_rotater1814_in[12], zll_main_rotater1814_in[24], zll_main_rotater1814_in[23], zll_main_rotater1814_in[22], zll_main_rotater1814_in[21], zll_main_rotater1814_in[20], zll_main_rotater1814_in[19], zll_main_rotater1814_in[18], zll_main_rotater1814_in[17], zll_main_rotater1814_in[16], zll_main_rotater1814_in[15], zll_main_rotater1814_in[14], zll_main_rotater1814_in[13], zll_main_rotater1814_in[11], zll_main_rotater1814_in[10], zll_main_rotater1814_in[9], zll_main_rotater1814_in[8], zll_main_rotater1814_in[7], zll_main_rotater1814_in[6], zll_main_rotater1814_in[5], zll_main_rotater1814_in[4], zll_main_rotater1814_in[3], zll_main_rotater1814_in[2], zll_main_rotater1814_in[1], zll_main_rotater1814_in[0]};
  assign zll_main_rotater184_in = {zll_main_rotater1815_in[31], zll_main_rotater1815_in[30], zll_main_rotater1815_in[29], zll_main_rotater1815_in[11], zll_main_rotater1815_in[28], zll_main_rotater1815_in[27], zll_main_rotater1815_in[26], zll_main_rotater1815_in[25], zll_main_rotater1815_in[24], zll_main_rotater1815_in[23], zll_main_rotater1815_in[22], zll_main_rotater1815_in[21], zll_main_rotater1815_in[20], zll_main_rotater1815_in[19], zll_main_rotater1815_in[18], zll_main_rotater1815_in[17], zll_main_rotater1815_in[16], zll_main_rotater1815_in[15], zll_main_rotater1815_in[14], zll_main_rotater1815_in[13], zll_main_rotater1815_in[12], zll_main_rotater1815_in[10], zll_main_rotater1815_in[9], zll_main_rotater1815_in[8], zll_main_rotater1815_in[7], zll_main_rotater1815_in[6], zll_main_rotater1815_in[5], zll_main_rotater1815_in[4], zll_main_rotater1815_in[3], zll_main_rotater1815_in[2], zll_main_rotater1815_in[1], zll_main_rotater1815_in[0]};
  assign zll_main_rotater182_in = {zll_main_rotater184_in[31], zll_main_rotater184_in[30], zll_main_rotater184_in[29], zll_main_rotater184_in[28], zll_main_rotater184_in[27], zll_main_rotater184_in[26], zll_main_rotater184_in[25], zll_main_rotater184_in[9], zll_main_rotater184_in[24], zll_main_rotater184_in[23], zll_main_rotater184_in[22], zll_main_rotater184_in[21], zll_main_rotater184_in[20], zll_main_rotater184_in[19], zll_main_rotater184_in[18], zll_main_rotater184_in[17], zll_main_rotater184_in[16], zll_main_rotater184_in[15], zll_main_rotater184_in[14], zll_main_rotater184_in[13], zll_main_rotater184_in[12], zll_main_rotater184_in[11], zll_main_rotater184_in[10], zll_main_rotater184_in[8], zll_main_rotater184_in[7], zll_main_rotater184_in[6], zll_main_rotater184_in[5], zll_main_rotater184_in[4], zll_main_rotater184_in[3], zll_main_rotater184_in[2], zll_main_rotater184_in[1], zll_main_rotater184_in[0]};
  assign zll_main_rotater1823_in = {zll_main_rotater182_in[31], zll_main_rotater182_in[30], zll_main_rotater182_in[29], zll_main_rotater182_in[28], zll_main_rotater182_in[27], zll_main_rotater182_in[26], zll_main_rotater182_in[25], zll_main_rotater182_in[24], zll_main_rotater182_in[8], zll_main_rotater182_in[23], zll_main_rotater182_in[22], zll_main_rotater182_in[21], zll_main_rotater182_in[20], zll_main_rotater182_in[19], zll_main_rotater182_in[18], zll_main_rotater182_in[17], zll_main_rotater182_in[16], zll_main_rotater182_in[15], zll_main_rotater182_in[14], zll_main_rotater182_in[13], zll_main_rotater182_in[12], zll_main_rotater182_in[11], zll_main_rotater182_in[10], zll_main_rotater182_in[9], zll_main_rotater182_in[7], zll_main_rotater182_in[6], zll_main_rotater182_in[5], zll_main_rotater182_in[4], zll_main_rotater182_in[3], zll_main_rotater182_in[2], zll_main_rotater182_in[1], zll_main_rotater182_in[0]};
  assign zll_main_rotater1829_in = {zll_main_rotater1823_in[31], zll_main_rotater1823_in[30], zll_main_rotater1823_in[29], zll_main_rotater1823_in[28], zll_main_rotater1823_in[27], zll_main_rotater1823_in[26], zll_main_rotater1823_in[25], zll_main_rotater1823_in[24], zll_main_rotater1823_in[23], zll_main_rotater1823_in[22], zll_main_rotater1823_in[21], zll_main_rotater1823_in[20], zll_main_rotater1823_in[19], zll_main_rotater1823_in[18], zll_main_rotater1823_in[17], zll_main_rotater1823_in[16], zll_main_rotater1823_in[15], zll_main_rotater1823_in[14], zll_main_rotater1823_in[13], zll_main_rotater1823_in[7], zll_main_rotater1823_in[12], zll_main_rotater1823_in[11], zll_main_rotater1823_in[10], zll_main_rotater1823_in[9], zll_main_rotater1823_in[8], zll_main_rotater1823_in[6], zll_main_rotater1823_in[5], zll_main_rotater1823_in[4], zll_main_rotater1823_in[3], zll_main_rotater1823_in[2], zll_main_rotater1823_in[1], zll_main_rotater1823_in[0]};
  assign zll_main_rotater1810_in = {zll_main_rotater1829_in[31], zll_main_rotater1829_in[30], zll_main_rotater1829_in[29], zll_main_rotater1829_in[28], zll_main_rotater1829_in[27], zll_main_rotater1829_in[26], zll_main_rotater1829_in[6], zll_main_rotater1829_in[25], zll_main_rotater1829_in[24], zll_main_rotater1829_in[23], zll_main_rotater1829_in[22], zll_main_rotater1829_in[21], zll_main_rotater1829_in[20], zll_main_rotater1829_in[19], zll_main_rotater1829_in[18], zll_main_rotater1829_in[17], zll_main_rotater1829_in[16], zll_main_rotater1829_in[15], zll_main_rotater1829_in[14], zll_main_rotater1829_in[13], zll_main_rotater1829_in[12], zll_main_rotater1829_in[11], zll_main_rotater1829_in[10], zll_main_rotater1829_in[9], zll_main_rotater1829_in[8], zll_main_rotater1829_in[7], zll_main_rotater1829_in[5], zll_main_rotater1829_in[4], zll_main_rotater1829_in[3], zll_main_rotater1829_in[2], zll_main_rotater1829_in[1], zll_main_rotater1829_in[0]};
  assign zll_main_rotater183_in = {zll_main_rotater1810_in[31], zll_main_rotater1810_in[30], zll_main_rotater1810_in[29], zll_main_rotater1810_in[28], zll_main_rotater1810_in[27], zll_main_rotater1810_in[26], zll_main_rotater1810_in[25], zll_main_rotater1810_in[24], zll_main_rotater1810_in[23], zll_main_rotater1810_in[22], zll_main_rotater1810_in[21], zll_main_rotater1810_in[20], zll_main_rotater1810_in[19], zll_main_rotater1810_in[18], zll_main_rotater1810_in[17], zll_main_rotater1810_in[16], zll_main_rotater1810_in[15], zll_main_rotater1810_in[14], zll_main_rotater1810_in[13], zll_main_rotater1810_in[12], zll_main_rotater1810_in[11], zll_main_rotater1810_in[10], zll_main_rotater1810_in[9], zll_main_rotater1810_in[5], zll_main_rotater1810_in[8], zll_main_rotater1810_in[7], zll_main_rotater1810_in[6], zll_main_rotater1810_in[4], zll_main_rotater1810_in[3], zll_main_rotater1810_in[2], zll_main_rotater1810_in[1], zll_main_rotater1810_in[0]};
  assign zll_main_rotater1816_in = {zll_main_rotater183_in[31], zll_main_rotater183_in[30], zll_main_rotater183_in[29], zll_main_rotater183_in[28], zll_main_rotater183_in[27], zll_main_rotater183_in[26], zll_main_rotater183_in[25], zll_main_rotater183_in[24], zll_main_rotater183_in[23], zll_main_rotater183_in[22], zll_main_rotater183_in[21], zll_main_rotater183_in[20], zll_main_rotater183_in[19], zll_main_rotater183_in[18], zll_main_rotater183_in[17], zll_main_rotater183_in[4], zll_main_rotater183_in[16], zll_main_rotater183_in[15], zll_main_rotater183_in[14], zll_main_rotater183_in[13], zll_main_rotater183_in[12], zll_main_rotater183_in[11], zll_main_rotater183_in[10], zll_main_rotater183_in[9], zll_main_rotater183_in[8], zll_main_rotater183_in[7], zll_main_rotater183_in[6], zll_main_rotater183_in[5], zll_main_rotater183_in[3], zll_main_rotater183_in[2], zll_main_rotater183_in[1], zll_main_rotater183_in[0]};
  assign zll_main_rotater189_in = {zll_main_rotater1816_in[31], zll_main_rotater1816_in[30], zll_main_rotater1816_in[3], zll_main_rotater1816_in[29], zll_main_rotater1816_in[28], zll_main_rotater1816_in[27], zll_main_rotater1816_in[26], zll_main_rotater1816_in[25], zll_main_rotater1816_in[24], zll_main_rotater1816_in[23], zll_main_rotater1816_in[22], zll_main_rotater1816_in[21], zll_main_rotater1816_in[20], zll_main_rotater1816_in[19], zll_main_rotater1816_in[18], zll_main_rotater1816_in[17], zll_main_rotater1816_in[16], zll_main_rotater1816_in[15], zll_main_rotater1816_in[14], zll_main_rotater1816_in[13], zll_main_rotater1816_in[12], zll_main_rotater1816_in[11], zll_main_rotater1816_in[10], zll_main_rotater1816_in[9], zll_main_rotater1816_in[8], zll_main_rotater1816_in[7], zll_main_rotater1816_in[6], zll_main_rotater1816_in[5], zll_main_rotater1816_in[4], zll_main_rotater1816_in[2], zll_main_rotater1816_in[1], zll_main_rotater1816_in[0]};
  assign zll_main_rotater18_in = {zll_main_rotater189_in[31], zll_main_rotater189_in[30], zll_main_rotater189_in[29], zll_main_rotater189_in[28], zll_main_rotater189_in[2], zll_main_rotater189_in[27], zll_main_rotater189_in[26], zll_main_rotater189_in[25], zll_main_rotater189_in[24], zll_main_rotater189_in[23], zll_main_rotater189_in[22], zll_main_rotater189_in[21], zll_main_rotater189_in[20], zll_main_rotater189_in[19], zll_main_rotater189_in[18], zll_main_rotater189_in[17], zll_main_rotater189_in[16], zll_main_rotater189_in[15], zll_main_rotater189_in[14], zll_main_rotater189_in[13], zll_main_rotater189_in[12], zll_main_rotater189_in[11], zll_main_rotater189_in[10], zll_main_rotater189_in[9], zll_main_rotater189_in[8], zll_main_rotater189_in[7], zll_main_rotater189_in[6], zll_main_rotater189_in[5], zll_main_rotater189_in[4], zll_main_rotater189_in[3], zll_main_rotater189_in[1], zll_main_rotater189_in[0]};
  assign zll_main_rotater1812_in = {zll_main_rotater18_in[31], zll_main_rotater18_in[30], zll_main_rotater18_in[29], zll_main_rotater18_in[28], zll_main_rotater18_in[27], zll_main_rotater18_in[26], zll_main_rotater18_in[25], zll_main_rotater18_in[24], zll_main_rotater18_in[23], zll_main_rotater18_in[22], zll_main_rotater18_in[21], zll_main_rotater18_in[1], zll_main_rotater18_in[20], zll_main_rotater18_in[19], zll_main_rotater18_in[18], zll_main_rotater18_in[17], zll_main_rotater18_in[16], zll_main_rotater18_in[15], zll_main_rotater18_in[14], zll_main_rotater18_in[13], zll_main_rotater18_in[12], zll_main_rotater18_in[11], zll_main_rotater18_in[10], zll_main_rotater18_in[9], zll_main_rotater18_in[8], zll_main_rotater18_in[7], zll_main_rotater18_in[6], zll_main_rotater18_in[5], zll_main_rotater18_in[4], zll_main_rotater18_in[3], zll_main_rotater18_in[2], zll_main_rotater18_in[0]};
  assign xorw32_inR2 = {{zll_main_rotater715_in[10], zll_main_rotater715_in[25], zll_main_rotater715_in[12], zll_main_rotater715_in[26], zll_main_rotater715_in[2], zll_main_rotater715_in[23], zll_main_rotater715_in[0], zll_main_rotater715_in[31], zll_main_rotater715_in[6], zll_main_rotater715_in[1], zll_main_rotater715_in[27], zll_main_rotater715_in[13], zll_main_rotater715_in[28], zll_main_rotater715_in[7], zll_main_rotater715_in[9], zll_main_rotater715_in[19], zll_main_rotater715_in[8], zll_main_rotater715_in[21], zll_main_rotater715_in[22], zll_main_rotater715_in[18], zll_main_rotater715_in[30], zll_main_rotater715_in[15], zll_main_rotater715_in[24], zll_main_rotater715_in[16], zll_main_rotater715_in[29], zll_main_rotater715_in[3], zll_main_rotater715_in[4], zll_main_rotater715_in[14], zll_main_rotater715_in[5], zll_main_rotater715_in[20], zll_main_rotater715_in[17], zll_main_rotater715_in[11]}, {zll_main_rotater1812_in[16], zll_main_rotater1812_in[28], zll_main_rotater1812_in[9], zll_main_rotater1812_in[25], zll_main_rotater1812_in[8], zll_main_rotater1812_in[17], zll_main_rotater1812_in[26], zll_main_rotater1812_in[1], zll_main_rotater1812_in[21], zll_main_rotater1812_in[19], zll_main_rotater1812_in[7], zll_main_rotater1812_in[23], zll_main_rotater1812_in[4], zll_main_rotater1812_in[13], zll_main_rotater1812_in[29], zll_main_rotater1812_in[27], zll_main_rotater1812_in[20], zll_main_rotater1812_in[0], zll_main_rotater1812_in[3], zll_main_rotater1812_in[14], zll_main_rotater1812_in[15], zll_main_rotater1812_in[11], zll_main_rotater1812_in[18], zll_main_rotater1812_in[30], zll_main_rotater1812_in[2], zll_main_rotater1812_in[22], zll_main_rotater1812_in[10], zll_main_rotater1812_in[24], zll_main_rotater1812_in[31], zll_main_rotater1812_in[5], zll_main_rotater1812_in[12], zll_main_rotater1812_in[6]}};
  xorW32  instR3 (xorw32_inR2[63:32], xorw32_inR2[31:0], extresR3[31:0]);
  assign main_shiftr3_in = main_sigma0_in[31:0];
  assign zll_main_shiftr311_in = main_shiftr3_in[31:0];
  assign zll_main_shiftr38_in = {zll_main_shiftr311_in[30], zll_main_shiftr311_in[31], zll_main_shiftr311_in[29], zll_main_shiftr311_in[28], zll_main_shiftr311_in[27], zll_main_shiftr311_in[26], zll_main_shiftr311_in[25], zll_main_shiftr311_in[24], zll_main_shiftr311_in[23], zll_main_shiftr311_in[22], zll_main_shiftr311_in[21], zll_main_shiftr311_in[20], zll_main_shiftr311_in[19], zll_main_shiftr311_in[18], zll_main_shiftr311_in[17], zll_main_shiftr311_in[16], zll_main_shiftr311_in[15], zll_main_shiftr311_in[14], zll_main_shiftr311_in[13], zll_main_shiftr311_in[12], zll_main_shiftr311_in[11], zll_main_shiftr311_in[10], zll_main_shiftr311_in[9], zll_main_shiftr311_in[8], zll_main_shiftr311_in[7], zll_main_shiftr311_in[6], zll_main_shiftr311_in[5], zll_main_shiftr311_in[4], zll_main_shiftr311_in[3], zll_main_shiftr311_in[2], zll_main_shiftr311_in[1], zll_main_shiftr311_in[0]};
  assign zll_main_shiftr330_in = {zll_main_shiftr38_in[31], zll_main_shiftr38_in[29], zll_main_shiftr38_in[30], zll_main_shiftr38_in[28], zll_main_shiftr38_in[27], zll_main_shiftr38_in[26], zll_main_shiftr38_in[25], zll_main_shiftr38_in[24], zll_main_shiftr38_in[23], zll_main_shiftr38_in[22], zll_main_shiftr38_in[21], zll_main_shiftr38_in[20], zll_main_shiftr38_in[19], zll_main_shiftr38_in[18], zll_main_shiftr38_in[17], zll_main_shiftr38_in[16], zll_main_shiftr38_in[15], zll_main_shiftr38_in[14], zll_main_shiftr38_in[13], zll_main_shiftr38_in[12], zll_main_shiftr38_in[11], zll_main_shiftr38_in[10], zll_main_shiftr38_in[9], zll_main_shiftr38_in[8], zll_main_shiftr38_in[7], zll_main_shiftr38_in[6], zll_main_shiftr38_in[5], zll_main_shiftr38_in[4], zll_main_shiftr38_in[3], zll_main_shiftr38_in[2], zll_main_shiftr38_in[1], zll_main_shiftr38_in[0]};
  assign zll_main_shiftr36_in = {zll_main_shiftr330_in[31], zll_main_shiftr330_in[27], zll_main_shiftr330_in[30], zll_main_shiftr330_in[29], zll_main_shiftr330_in[28], zll_main_shiftr330_in[26], zll_main_shiftr330_in[25], zll_main_shiftr330_in[24], zll_main_shiftr330_in[23], zll_main_shiftr330_in[22], zll_main_shiftr330_in[21], zll_main_shiftr330_in[20], zll_main_shiftr330_in[19], zll_main_shiftr330_in[18], zll_main_shiftr330_in[17], zll_main_shiftr330_in[16], zll_main_shiftr330_in[15], zll_main_shiftr330_in[14], zll_main_shiftr330_in[13], zll_main_shiftr330_in[12], zll_main_shiftr330_in[11], zll_main_shiftr330_in[10], zll_main_shiftr330_in[9], zll_main_shiftr330_in[8], zll_main_shiftr330_in[7], zll_main_shiftr330_in[6], zll_main_shiftr330_in[5], zll_main_shiftr330_in[4], zll_main_shiftr330_in[3], zll_main_shiftr330_in[2], zll_main_shiftr330_in[1], zll_main_shiftr330_in[0]};
  assign zll_main_shiftr312_in = {zll_main_shiftr36_in[31], zll_main_shiftr36_in[30], zll_main_shiftr36_in[29], zll_main_shiftr36_in[25], zll_main_shiftr36_in[28], zll_main_shiftr36_in[27], zll_main_shiftr36_in[26], zll_main_shiftr36_in[24], zll_main_shiftr36_in[23], zll_main_shiftr36_in[22], zll_main_shiftr36_in[21], zll_main_shiftr36_in[20], zll_main_shiftr36_in[19], zll_main_shiftr36_in[18], zll_main_shiftr36_in[17], zll_main_shiftr36_in[16], zll_main_shiftr36_in[15], zll_main_shiftr36_in[14], zll_main_shiftr36_in[13], zll_main_shiftr36_in[12], zll_main_shiftr36_in[11], zll_main_shiftr36_in[10], zll_main_shiftr36_in[9], zll_main_shiftr36_in[8], zll_main_shiftr36_in[7], zll_main_shiftr36_in[6], zll_main_shiftr36_in[5], zll_main_shiftr36_in[4], zll_main_shiftr36_in[3], zll_main_shiftr36_in[2], zll_main_shiftr36_in[1], zll_main_shiftr36_in[0]};
  assign zll_main_shiftr326_in = {zll_main_shiftr312_in[31], zll_main_shiftr312_in[24], zll_main_shiftr312_in[30], zll_main_shiftr312_in[29], zll_main_shiftr312_in[28], zll_main_shiftr312_in[27], zll_main_shiftr312_in[26], zll_main_shiftr312_in[25], zll_main_shiftr312_in[23], zll_main_shiftr312_in[22], zll_main_shiftr312_in[21], zll_main_shiftr312_in[20], zll_main_shiftr312_in[19], zll_main_shiftr312_in[18], zll_main_shiftr312_in[17], zll_main_shiftr312_in[16], zll_main_shiftr312_in[15], zll_main_shiftr312_in[14], zll_main_shiftr312_in[13], zll_main_shiftr312_in[12], zll_main_shiftr312_in[11], zll_main_shiftr312_in[10], zll_main_shiftr312_in[9], zll_main_shiftr312_in[8], zll_main_shiftr312_in[7], zll_main_shiftr312_in[6], zll_main_shiftr312_in[5], zll_main_shiftr312_in[4], zll_main_shiftr312_in[3], zll_main_shiftr312_in[2], zll_main_shiftr312_in[1], zll_main_shiftr312_in[0]};
  assign zll_main_shiftr322_in = {zll_main_shiftr326_in[31], zll_main_shiftr326_in[30], zll_main_shiftr326_in[23], zll_main_shiftr326_in[29], zll_main_shiftr326_in[28], zll_main_shiftr326_in[27], zll_main_shiftr326_in[26], zll_main_shiftr326_in[25], zll_main_shiftr326_in[24], zll_main_shiftr326_in[22], zll_main_shiftr326_in[21], zll_main_shiftr326_in[20], zll_main_shiftr326_in[19], zll_main_shiftr326_in[18], zll_main_shiftr326_in[17], zll_main_shiftr326_in[16], zll_main_shiftr326_in[15], zll_main_shiftr326_in[14], zll_main_shiftr326_in[13], zll_main_shiftr326_in[12], zll_main_shiftr326_in[11], zll_main_shiftr326_in[10], zll_main_shiftr326_in[9], zll_main_shiftr326_in[8], zll_main_shiftr326_in[7], zll_main_shiftr326_in[6], zll_main_shiftr326_in[5], zll_main_shiftr326_in[4], zll_main_shiftr326_in[3], zll_main_shiftr326_in[2], zll_main_shiftr326_in[1], zll_main_shiftr326_in[0]};
  assign zll_main_shiftr321_in = {zll_main_shiftr322_in[31], zll_main_shiftr322_in[30], zll_main_shiftr322_in[22], zll_main_shiftr322_in[29], zll_main_shiftr322_in[28], zll_main_shiftr322_in[27], zll_main_shiftr322_in[26], zll_main_shiftr322_in[25], zll_main_shiftr322_in[24], zll_main_shiftr322_in[23], zll_main_shiftr322_in[21], zll_main_shiftr322_in[20], zll_main_shiftr322_in[19], zll_main_shiftr322_in[18], zll_main_shiftr322_in[17], zll_main_shiftr322_in[16], zll_main_shiftr322_in[15], zll_main_shiftr322_in[14], zll_main_shiftr322_in[13], zll_main_shiftr322_in[12], zll_main_shiftr322_in[11], zll_main_shiftr322_in[10], zll_main_shiftr322_in[9], zll_main_shiftr322_in[8], zll_main_shiftr322_in[7], zll_main_shiftr322_in[6], zll_main_shiftr322_in[5], zll_main_shiftr322_in[4], zll_main_shiftr322_in[3], zll_main_shiftr322_in[2], zll_main_shiftr322_in[1], zll_main_shiftr322_in[0]};
  assign zll_main_shiftr316_in = {zll_main_shiftr321_in[21], zll_main_shiftr321_in[31], zll_main_shiftr321_in[30], zll_main_shiftr321_in[29], zll_main_shiftr321_in[28], zll_main_shiftr321_in[27], zll_main_shiftr321_in[26], zll_main_shiftr321_in[25], zll_main_shiftr321_in[24], zll_main_shiftr321_in[23], zll_main_shiftr321_in[22], zll_main_shiftr321_in[20], zll_main_shiftr321_in[19], zll_main_shiftr321_in[18], zll_main_shiftr321_in[17], zll_main_shiftr321_in[16], zll_main_shiftr321_in[15], zll_main_shiftr321_in[14], zll_main_shiftr321_in[13], zll_main_shiftr321_in[12], zll_main_shiftr321_in[11], zll_main_shiftr321_in[10], zll_main_shiftr321_in[9], zll_main_shiftr321_in[8], zll_main_shiftr321_in[7], zll_main_shiftr321_in[6], zll_main_shiftr321_in[5], zll_main_shiftr321_in[4], zll_main_shiftr321_in[3], zll_main_shiftr321_in[2], zll_main_shiftr321_in[1], zll_main_shiftr321_in[0]};
  assign zll_main_shiftr323_in = {zll_main_shiftr316_in[31], zll_main_shiftr316_in[30], zll_main_shiftr316_in[29], zll_main_shiftr316_in[20], zll_main_shiftr316_in[28], zll_main_shiftr316_in[27], zll_main_shiftr316_in[26], zll_main_shiftr316_in[25], zll_main_shiftr316_in[24], zll_main_shiftr316_in[23], zll_main_shiftr316_in[22], zll_main_shiftr316_in[21], zll_main_shiftr316_in[19], zll_main_shiftr316_in[18], zll_main_shiftr316_in[17], zll_main_shiftr316_in[16], zll_main_shiftr316_in[15], zll_main_shiftr316_in[14], zll_main_shiftr316_in[13], zll_main_shiftr316_in[12], zll_main_shiftr316_in[11], zll_main_shiftr316_in[10], zll_main_shiftr316_in[9], zll_main_shiftr316_in[8], zll_main_shiftr316_in[7], zll_main_shiftr316_in[6], zll_main_shiftr316_in[5], zll_main_shiftr316_in[4], zll_main_shiftr316_in[3], zll_main_shiftr316_in[2], zll_main_shiftr316_in[1], zll_main_shiftr316_in[0]};
  assign zll_main_shiftr3_in = {zll_main_shiftr323_in[31], zll_main_shiftr323_in[30], zll_main_shiftr323_in[29], zll_main_shiftr323_in[28], zll_main_shiftr323_in[27], zll_main_shiftr323_in[26], zll_main_shiftr323_in[25], zll_main_shiftr323_in[19], zll_main_shiftr323_in[24], zll_main_shiftr323_in[23], zll_main_shiftr323_in[22], zll_main_shiftr323_in[21], zll_main_shiftr323_in[20], zll_main_shiftr323_in[18], zll_main_shiftr323_in[17], zll_main_shiftr323_in[16], zll_main_shiftr323_in[15], zll_main_shiftr323_in[14], zll_main_shiftr323_in[13], zll_main_shiftr323_in[12], zll_main_shiftr323_in[11], zll_main_shiftr323_in[10], zll_main_shiftr323_in[9], zll_main_shiftr323_in[8], zll_main_shiftr323_in[7], zll_main_shiftr323_in[6], zll_main_shiftr323_in[5], zll_main_shiftr323_in[4], zll_main_shiftr323_in[3], zll_main_shiftr323_in[2], zll_main_shiftr323_in[1], zll_main_shiftr323_in[0]};
  assign zll_main_shiftr33_in = {zll_main_shiftr3_in[31], zll_main_shiftr3_in[30], zll_main_shiftr3_in[29], zll_main_shiftr3_in[28], zll_main_shiftr3_in[27], zll_main_shiftr3_in[26], zll_main_shiftr3_in[25], zll_main_shiftr3_in[24], zll_main_shiftr3_in[23], zll_main_shiftr3_in[22], zll_main_shiftr3_in[18], zll_main_shiftr3_in[21], zll_main_shiftr3_in[20], zll_main_shiftr3_in[19], zll_main_shiftr3_in[17], zll_main_shiftr3_in[16], zll_main_shiftr3_in[15], zll_main_shiftr3_in[14], zll_main_shiftr3_in[13], zll_main_shiftr3_in[12], zll_main_shiftr3_in[11], zll_main_shiftr3_in[10], zll_main_shiftr3_in[9], zll_main_shiftr3_in[8], zll_main_shiftr3_in[7], zll_main_shiftr3_in[6], zll_main_shiftr3_in[5], zll_main_shiftr3_in[4], zll_main_shiftr3_in[3], zll_main_shiftr3_in[2], zll_main_shiftr3_in[1], zll_main_shiftr3_in[0]};
  assign zll_main_shiftr310_in = {zll_main_shiftr33_in[31], zll_main_shiftr33_in[17], zll_main_shiftr33_in[30], zll_main_shiftr33_in[29], zll_main_shiftr33_in[28], zll_main_shiftr33_in[27], zll_main_shiftr33_in[26], zll_main_shiftr33_in[25], zll_main_shiftr33_in[24], zll_main_shiftr33_in[23], zll_main_shiftr33_in[22], zll_main_shiftr33_in[21], zll_main_shiftr33_in[20], zll_main_shiftr33_in[19], zll_main_shiftr33_in[18], zll_main_shiftr33_in[16], zll_main_shiftr33_in[15], zll_main_shiftr33_in[14], zll_main_shiftr33_in[13], zll_main_shiftr33_in[12], zll_main_shiftr33_in[11], zll_main_shiftr33_in[10], zll_main_shiftr33_in[9], zll_main_shiftr33_in[8], zll_main_shiftr33_in[7], zll_main_shiftr33_in[6], zll_main_shiftr33_in[5], zll_main_shiftr33_in[4], zll_main_shiftr33_in[3], zll_main_shiftr33_in[2], zll_main_shiftr33_in[1], zll_main_shiftr33_in[0]};
  assign zll_main_shiftr39_in = {zll_main_shiftr310_in[31], zll_main_shiftr310_in[30], zll_main_shiftr310_in[29], zll_main_shiftr310_in[28], zll_main_shiftr310_in[27], zll_main_shiftr310_in[26], zll_main_shiftr310_in[25], zll_main_shiftr310_in[24], zll_main_shiftr310_in[23], zll_main_shiftr310_in[22], zll_main_shiftr310_in[21], zll_main_shiftr310_in[20], zll_main_shiftr310_in[16], zll_main_shiftr310_in[19], zll_main_shiftr310_in[18], zll_main_shiftr310_in[17], zll_main_shiftr310_in[15], zll_main_shiftr310_in[14], zll_main_shiftr310_in[13], zll_main_shiftr310_in[12], zll_main_shiftr310_in[11], zll_main_shiftr310_in[10], zll_main_shiftr310_in[9], zll_main_shiftr310_in[8], zll_main_shiftr310_in[7], zll_main_shiftr310_in[6], zll_main_shiftr310_in[5], zll_main_shiftr310_in[4], zll_main_shiftr310_in[3], zll_main_shiftr310_in[2], zll_main_shiftr310_in[1], zll_main_shiftr310_in[0]};
  assign zll_main_shiftr320_in = {zll_main_shiftr39_in[31], zll_main_shiftr39_in[30], zll_main_shiftr39_in[29], zll_main_shiftr39_in[28], zll_main_shiftr39_in[27], zll_main_shiftr39_in[26], zll_main_shiftr39_in[25], zll_main_shiftr39_in[24], zll_main_shiftr39_in[23], zll_main_shiftr39_in[22], zll_main_shiftr39_in[21], zll_main_shiftr39_in[20], zll_main_shiftr39_in[19], zll_main_shiftr39_in[18], zll_main_shiftr39_in[15], zll_main_shiftr39_in[17], zll_main_shiftr39_in[16], zll_main_shiftr39_in[14], zll_main_shiftr39_in[13], zll_main_shiftr39_in[12], zll_main_shiftr39_in[11], zll_main_shiftr39_in[10], zll_main_shiftr39_in[9], zll_main_shiftr39_in[8], zll_main_shiftr39_in[7], zll_main_shiftr39_in[6], zll_main_shiftr39_in[5], zll_main_shiftr39_in[4], zll_main_shiftr39_in[3], zll_main_shiftr39_in[2], zll_main_shiftr39_in[1], zll_main_shiftr39_in[0]};
  assign zll_main_shiftr327_in = {zll_main_shiftr320_in[31], zll_main_shiftr320_in[30], zll_main_shiftr320_in[29], zll_main_shiftr320_in[28], zll_main_shiftr320_in[27], zll_main_shiftr320_in[26], zll_main_shiftr320_in[25], zll_main_shiftr320_in[24], zll_main_shiftr320_in[14], zll_main_shiftr320_in[23], zll_main_shiftr320_in[22], zll_main_shiftr320_in[21], zll_main_shiftr320_in[20], zll_main_shiftr320_in[19], zll_main_shiftr320_in[18], zll_main_shiftr320_in[17], zll_main_shiftr320_in[16], zll_main_shiftr320_in[15], zll_main_shiftr320_in[13], zll_main_shiftr320_in[12], zll_main_shiftr320_in[11], zll_main_shiftr320_in[10], zll_main_shiftr320_in[9], zll_main_shiftr320_in[8], zll_main_shiftr320_in[7], zll_main_shiftr320_in[6], zll_main_shiftr320_in[5], zll_main_shiftr320_in[4], zll_main_shiftr320_in[3], zll_main_shiftr320_in[2], zll_main_shiftr320_in[1], zll_main_shiftr320_in[0]};
  assign zll_main_shiftr315_in = {zll_main_shiftr327_in[31], zll_main_shiftr327_in[30], zll_main_shiftr327_in[29], zll_main_shiftr327_in[28], zll_main_shiftr327_in[27], zll_main_shiftr327_in[26], zll_main_shiftr327_in[13], zll_main_shiftr327_in[25], zll_main_shiftr327_in[24], zll_main_shiftr327_in[23], zll_main_shiftr327_in[22], zll_main_shiftr327_in[21], zll_main_shiftr327_in[20], zll_main_shiftr327_in[19], zll_main_shiftr327_in[18], zll_main_shiftr327_in[17], zll_main_shiftr327_in[16], zll_main_shiftr327_in[15], zll_main_shiftr327_in[14], zll_main_shiftr327_in[12], zll_main_shiftr327_in[11], zll_main_shiftr327_in[10], zll_main_shiftr327_in[9], zll_main_shiftr327_in[8], zll_main_shiftr327_in[7], zll_main_shiftr327_in[6], zll_main_shiftr327_in[5], zll_main_shiftr327_in[4], zll_main_shiftr327_in[3], zll_main_shiftr327_in[2], zll_main_shiftr327_in[1], zll_main_shiftr327_in[0]};
  assign zll_main_shiftr329_in = {zll_main_shiftr315_in[31], zll_main_shiftr315_in[30], zll_main_shiftr315_in[29], zll_main_shiftr315_in[28], zll_main_shiftr315_in[27], zll_main_shiftr315_in[12], zll_main_shiftr315_in[26], zll_main_shiftr315_in[25], zll_main_shiftr315_in[24], zll_main_shiftr315_in[23], zll_main_shiftr315_in[22], zll_main_shiftr315_in[21], zll_main_shiftr315_in[20], zll_main_shiftr315_in[19], zll_main_shiftr315_in[18], zll_main_shiftr315_in[17], zll_main_shiftr315_in[16], zll_main_shiftr315_in[15], zll_main_shiftr315_in[14], zll_main_shiftr315_in[13], zll_main_shiftr315_in[11], zll_main_shiftr315_in[10], zll_main_shiftr315_in[9], zll_main_shiftr315_in[8], zll_main_shiftr315_in[7], zll_main_shiftr315_in[6], zll_main_shiftr315_in[5], zll_main_shiftr315_in[4], zll_main_shiftr315_in[3], zll_main_shiftr315_in[2], zll_main_shiftr315_in[1], zll_main_shiftr315_in[0]};
  assign zll_main_shiftr331_in = {zll_main_shiftr329_in[31], zll_main_shiftr329_in[11], zll_main_shiftr329_in[30], zll_main_shiftr329_in[29], zll_main_shiftr329_in[28], zll_main_shiftr329_in[27], zll_main_shiftr329_in[26], zll_main_shiftr329_in[25], zll_main_shiftr329_in[24], zll_main_shiftr329_in[23], zll_main_shiftr329_in[22], zll_main_shiftr329_in[21], zll_main_shiftr329_in[20], zll_main_shiftr329_in[19], zll_main_shiftr329_in[18], zll_main_shiftr329_in[17], zll_main_shiftr329_in[16], zll_main_shiftr329_in[15], zll_main_shiftr329_in[14], zll_main_shiftr329_in[13], zll_main_shiftr329_in[12], zll_main_shiftr329_in[10], zll_main_shiftr329_in[9], zll_main_shiftr329_in[8], zll_main_shiftr329_in[7], zll_main_shiftr329_in[6], zll_main_shiftr329_in[5], zll_main_shiftr329_in[4], zll_main_shiftr329_in[3], zll_main_shiftr329_in[2], zll_main_shiftr329_in[1], zll_main_shiftr329_in[0]};
  assign zll_main_shiftr324_in = {zll_main_shiftr331_in[10], zll_main_shiftr331_in[31], zll_main_shiftr331_in[30], zll_main_shiftr331_in[29], zll_main_shiftr331_in[28], zll_main_shiftr331_in[27], zll_main_shiftr331_in[26], zll_main_shiftr331_in[25], zll_main_shiftr331_in[24], zll_main_shiftr331_in[23], zll_main_shiftr331_in[22], zll_main_shiftr331_in[21], zll_main_shiftr331_in[20], zll_main_shiftr331_in[19], zll_main_shiftr331_in[18], zll_main_shiftr331_in[17], zll_main_shiftr331_in[16], zll_main_shiftr331_in[15], zll_main_shiftr331_in[14], zll_main_shiftr331_in[13], zll_main_shiftr331_in[12], zll_main_shiftr331_in[11], zll_main_shiftr331_in[9], zll_main_shiftr331_in[8], zll_main_shiftr331_in[7], zll_main_shiftr331_in[6], zll_main_shiftr331_in[5], zll_main_shiftr331_in[4], zll_main_shiftr331_in[3], zll_main_shiftr331_in[2], zll_main_shiftr331_in[1], zll_main_shiftr331_in[0]};
  assign zll_main_shiftr32_in = {zll_main_shiftr324_in[31], zll_main_shiftr324_in[30], zll_main_shiftr324_in[29], zll_main_shiftr324_in[28], zll_main_shiftr324_in[9], zll_main_shiftr324_in[27], zll_main_shiftr324_in[26], zll_main_shiftr324_in[25], zll_main_shiftr324_in[24], zll_main_shiftr324_in[23], zll_main_shiftr324_in[22], zll_main_shiftr324_in[21], zll_main_shiftr324_in[20], zll_main_shiftr324_in[19], zll_main_shiftr324_in[18], zll_main_shiftr324_in[17], zll_main_shiftr324_in[16], zll_main_shiftr324_in[15], zll_main_shiftr324_in[14], zll_main_shiftr324_in[13], zll_main_shiftr324_in[12], zll_main_shiftr324_in[11], zll_main_shiftr324_in[10], zll_main_shiftr324_in[8], zll_main_shiftr324_in[7], zll_main_shiftr324_in[6], zll_main_shiftr324_in[5], zll_main_shiftr324_in[4], zll_main_shiftr324_in[3], zll_main_shiftr324_in[2], zll_main_shiftr324_in[1], zll_main_shiftr324_in[0]};
  assign zll_main_shiftr325_in = {zll_main_shiftr32_in[31], zll_main_shiftr32_in[30], zll_main_shiftr32_in[29], zll_main_shiftr32_in[28], zll_main_shiftr32_in[27], zll_main_shiftr32_in[26], zll_main_shiftr32_in[25], zll_main_shiftr32_in[24], zll_main_shiftr32_in[23], zll_main_shiftr32_in[22], zll_main_shiftr32_in[21], zll_main_shiftr32_in[20], zll_main_shiftr32_in[19], zll_main_shiftr32_in[18], zll_main_shiftr32_in[17], zll_main_shiftr32_in[16], zll_main_shiftr32_in[15], zll_main_shiftr32_in[14], zll_main_shiftr32_in[13], zll_main_shiftr32_in[8], zll_main_shiftr32_in[12], zll_main_shiftr32_in[11], zll_main_shiftr32_in[10], zll_main_shiftr32_in[9], zll_main_shiftr32_in[7], zll_main_shiftr32_in[6], zll_main_shiftr32_in[5], zll_main_shiftr32_in[4], zll_main_shiftr32_in[3], zll_main_shiftr32_in[2], zll_main_shiftr32_in[1], zll_main_shiftr32_in[0]};
  assign zll_main_shiftr314_in = {zll_main_shiftr325_in[7], zll_main_shiftr325_in[31], zll_main_shiftr325_in[30], zll_main_shiftr325_in[29], zll_main_shiftr325_in[28], zll_main_shiftr325_in[27], zll_main_shiftr325_in[26], zll_main_shiftr325_in[25], zll_main_shiftr325_in[24], zll_main_shiftr325_in[23], zll_main_shiftr325_in[22], zll_main_shiftr325_in[21], zll_main_shiftr325_in[20], zll_main_shiftr325_in[19], zll_main_shiftr325_in[18], zll_main_shiftr325_in[17], zll_main_shiftr325_in[16], zll_main_shiftr325_in[15], zll_main_shiftr325_in[14], zll_main_shiftr325_in[13], zll_main_shiftr325_in[12], zll_main_shiftr325_in[11], zll_main_shiftr325_in[10], zll_main_shiftr325_in[9], zll_main_shiftr325_in[8], zll_main_shiftr325_in[6], zll_main_shiftr325_in[5], zll_main_shiftr325_in[4], zll_main_shiftr325_in[3], zll_main_shiftr325_in[2], zll_main_shiftr325_in[1], zll_main_shiftr325_in[0]};
  assign zll_main_shiftr35_in = {zll_main_shiftr314_in[31], zll_main_shiftr314_in[30], zll_main_shiftr314_in[29], zll_main_shiftr314_in[28], zll_main_shiftr314_in[27], zll_main_shiftr314_in[26], zll_main_shiftr314_in[25], zll_main_shiftr314_in[24], zll_main_shiftr314_in[23], zll_main_shiftr314_in[22], zll_main_shiftr314_in[21], zll_main_shiftr314_in[20], zll_main_shiftr314_in[19], zll_main_shiftr314_in[18], zll_main_shiftr314_in[17], zll_main_shiftr314_in[16], zll_main_shiftr314_in[15], zll_main_shiftr314_in[14], zll_main_shiftr314_in[13], zll_main_shiftr314_in[12], zll_main_shiftr314_in[11], zll_main_shiftr314_in[10], zll_main_shiftr314_in[9], zll_main_shiftr314_in[6], zll_main_shiftr314_in[8], zll_main_shiftr314_in[7], zll_main_shiftr314_in[5], zll_main_shiftr314_in[4], zll_main_shiftr314_in[3], zll_main_shiftr314_in[2], zll_main_shiftr314_in[1], zll_main_shiftr314_in[0]};
  assign zll_main_shiftr31_in = {zll_main_shiftr35_in[31], zll_main_shiftr35_in[5], zll_main_shiftr35_in[30], zll_main_shiftr35_in[29], zll_main_shiftr35_in[28], zll_main_shiftr35_in[27], zll_main_shiftr35_in[26], zll_main_shiftr35_in[25], zll_main_shiftr35_in[24], zll_main_shiftr35_in[23], zll_main_shiftr35_in[22], zll_main_shiftr35_in[21], zll_main_shiftr35_in[20], zll_main_shiftr35_in[19], zll_main_shiftr35_in[18], zll_main_shiftr35_in[17], zll_main_shiftr35_in[16], zll_main_shiftr35_in[15], zll_main_shiftr35_in[14], zll_main_shiftr35_in[13], zll_main_shiftr35_in[12], zll_main_shiftr35_in[11], zll_main_shiftr35_in[10], zll_main_shiftr35_in[9], zll_main_shiftr35_in[8], zll_main_shiftr35_in[7], zll_main_shiftr35_in[6], zll_main_shiftr35_in[4], zll_main_shiftr35_in[3], zll_main_shiftr35_in[2], zll_main_shiftr35_in[1], zll_main_shiftr35_in[0]};
  assign zll_main_shiftr37_in = {zll_main_shiftr31_in[31], zll_main_shiftr31_in[30], zll_main_shiftr31_in[29], zll_main_shiftr31_in[28], zll_main_shiftr31_in[27], zll_main_shiftr31_in[4], zll_main_shiftr31_in[26], zll_main_shiftr31_in[25], zll_main_shiftr31_in[24], zll_main_shiftr31_in[23], zll_main_shiftr31_in[22], zll_main_shiftr31_in[21], zll_main_shiftr31_in[20], zll_main_shiftr31_in[19], zll_main_shiftr31_in[18], zll_main_shiftr31_in[17], zll_main_shiftr31_in[16], zll_main_shiftr31_in[15], zll_main_shiftr31_in[14], zll_main_shiftr31_in[13], zll_main_shiftr31_in[12], zll_main_shiftr31_in[11], zll_main_shiftr31_in[10], zll_main_shiftr31_in[9], zll_main_shiftr31_in[8], zll_main_shiftr31_in[7], zll_main_shiftr31_in[6], zll_main_shiftr31_in[5], zll_main_shiftr31_in[3], zll_main_shiftr31_in[2], zll_main_shiftr31_in[1], zll_main_shiftr31_in[0]};
  assign zll_main_shiftr313_in = {zll_main_shiftr37_in[31], zll_main_shiftr37_in[30], zll_main_shiftr37_in[29], zll_main_shiftr37_in[28], zll_main_shiftr37_in[27], zll_main_shiftr37_in[26], zll_main_shiftr37_in[25], zll_main_shiftr37_in[24], zll_main_shiftr37_in[23], zll_main_shiftr37_in[22], zll_main_shiftr37_in[21], zll_main_shiftr37_in[20], zll_main_shiftr37_in[19], zll_main_shiftr37_in[18], zll_main_shiftr37_in[17], zll_main_shiftr37_in[16], zll_main_shiftr37_in[15], zll_main_shiftr37_in[14], zll_main_shiftr37_in[13], zll_main_shiftr37_in[12], zll_main_shiftr37_in[11], zll_main_shiftr37_in[10], zll_main_shiftr37_in[9], zll_main_shiftr37_in[8], zll_main_shiftr37_in[7], zll_main_shiftr37_in[6], zll_main_shiftr37_in[5], zll_main_shiftr37_in[3], zll_main_shiftr37_in[4], zll_main_shiftr37_in[2], zll_main_shiftr37_in[1], zll_main_shiftr37_in[0]};
  assign zll_main_shiftr328_in = {zll_main_shiftr313_in[31], zll_main_shiftr313_in[30], zll_main_shiftr313_in[29], zll_main_shiftr313_in[28], zll_main_shiftr313_in[27], zll_main_shiftr313_in[26], zll_main_shiftr313_in[25], zll_main_shiftr313_in[24], zll_main_shiftr313_in[23], zll_main_shiftr313_in[22], zll_main_shiftr313_in[21], zll_main_shiftr313_in[20], zll_main_shiftr313_in[19], zll_main_shiftr313_in[18], zll_main_shiftr313_in[17], zll_main_shiftr313_in[16], zll_main_shiftr313_in[15], zll_main_shiftr313_in[14], zll_main_shiftr313_in[13], zll_main_shiftr313_in[12], zll_main_shiftr313_in[11], zll_main_shiftr313_in[10], zll_main_shiftr313_in[9], zll_main_shiftr313_in[8], zll_main_shiftr313_in[7], zll_main_shiftr313_in[6], zll_main_shiftr313_in[5], zll_main_shiftr313_in[4], zll_main_shiftr313_in[3], zll_main_shiftr313_in[1], zll_main_shiftr313_in[0]};
  assign zll_main_shiftr34_in = {zll_main_shiftr328_in[30], zll_main_shiftr328_in[29], zll_main_shiftr328_in[28], zll_main_shiftr328_in[27], zll_main_shiftr328_in[26], zll_main_shiftr328_in[25], zll_main_shiftr328_in[24], zll_main_shiftr328_in[23], zll_main_shiftr328_in[22], zll_main_shiftr328_in[21], zll_main_shiftr328_in[20], zll_main_shiftr328_in[19], zll_main_shiftr328_in[18], zll_main_shiftr328_in[17], zll_main_shiftr328_in[16], zll_main_shiftr328_in[15], zll_main_shiftr328_in[14], zll_main_shiftr328_in[13], zll_main_shiftr328_in[12], zll_main_shiftr328_in[11], zll_main_shiftr328_in[10], zll_main_shiftr328_in[9], zll_main_shiftr328_in[8], zll_main_shiftr328_in[7], zll_main_shiftr328_in[6], zll_main_shiftr328_in[5], zll_main_shiftr328_in[4], zll_main_shiftr328_in[3], zll_main_shiftr328_in[2], zll_main_shiftr328_in[0]};
  assign xorw32_inR3 = {extresR3, {3'h0, zll_main_shiftr34_in[6], zll_main_shiftr34_in[21], zll_main_shiftr34_in[11], zll_main_shiftr34_in[3], zll_main_shiftr34_in[14], zll_main_shiftr34_in[1], zll_main_shiftr34_in[10], zll_main_shiftr34_in[20], zll_main_shiftr34_in[15], zll_main_shiftr34_in[17], zll_main_shiftr34_in[26], zll_main_shiftr34_in[19], zll_main_shiftr34_in[12], zll_main_shiftr34_in[9], zll_main_shiftr34_in[23], zll_main_shiftr34_in[8], zll_main_shiftr34_in[5], zll_main_shiftr34_in[13], zll_main_shiftr34_in[16], zll_main_shiftr34_in[18], zll_main_shiftr34_in[25], zll_main_shiftr34_in[27], zll_main_shiftr34_in[22], zll_main_shiftr34_in[7], zll_main_shiftr34_in[29], zll_main_shiftr34_in[4], zll_main_shiftr34_in[28], zll_main_shiftr34_in[24], zll_main_shiftr34_in[2]}};
  xorW32  instR4 (xorw32_inR3[63:32], xorw32_inR3[31:0], extresR4[31:0]);
  assign plusw32_inR1 = {extresR4, zll_main_updatesched2_in[159:128]};
  plusW32  instR5 (plusw32_inR1[63:32], plusw32_inR1[31:0], extresR5[31:0]);
  assign plusw32_inR2 = {extresR2, extresR5};
  plusW32  instR6 (plusw32_inR2[63:32], plusw32_inR2[31:0], extresR6[31:0]);
  assign zll_main_loop74_in = {zll_main_loop141_in[1093:1062], zll_main_loop141_in[1029:774], {zll_main_updatesched2_in[383:352], zll_main_updatesched2_in[447:416], zll_main_updatesched2_in[319:288], zll_main_updatesched2_in[95:64], zll_main_updatesched2_in[287:256], zll_main_updatesched2_in[191:160], zll_main_updatesched2_in[479:448], zll_main_updatesched2_in[127:96], zll_main_updatesched2_in[415:384], zll_main_updatesched2_in[511:480], zll_main_updatesched2_in[223:192], zll_main_updatesched2_in[255:224], zll_main_updatesched2_in[351:320], zll_main_updatesched2_in[63:32], zll_main_updatesched2_in[31:0], extresR6}, zll_main_loop141_in[261:6], zll_main_loop141_in[5:0]};
  assign zll_main_loop58_in = {zll_main_loop74_in[1061:1030], zll_main_loop74_in[1029:0]};
  assign zll_main_loop17_in = {zll_main_loop58_in[1061:1030], zll_main_loop58_in[773:262], zll_main_loop58_in[1029:774], zll_main_loop58_in[261:6], zll_main_loop58_in[5:0]};
  assign zll_main_loop151_in = {zll_main_loop42_in[1035:1030], {zll_main_loop17_in[1061:1030], zll_main_loop17_in[517:262], zll_main_loop17_in[1029:518], zll_main_loop17_in[261:6], zll_main_loop17_in[5:0]}};
  assign zll_main_loop20_in = {zll_main_loop151_in[1067:1062], zll_main_loop151_in[1061:0]};
  assign zll_main_loop32_in = {zll_main_loop20_in[1029:774], zll_main_loop20_in[1067:1062], zll_main_loop20_in[1061:1030], zll_main_loop20_in[773:262], zll_main_loop20_in[261:6], zll_main_loop20_in[5:0]};
  assign zll_main_loop103_in = {zll_main_loop32_in[1067:812], zll_main_loop32_in[773:262], zll_main_loop32_in[811:806], zll_main_loop32_in[805:774], zll_main_loop32_in[261:6], zll_main_loop32_in[5:0]};
  assign zll_main_loop72_in = {zll_main_loop103_in[299:294], zll_main_loop103_in[293:262], zll_main_loop103_in[1067:812], zll_main_loop103_in[811:300], zll_main_loop103_in[261:6], zll_main_loop103_in[5:0]};
  assign zll_main_loop15_in = {zll_main_loop72_in[1061:1030], zll_main_loop72_in[1067:1062], zll_main_loop72_in[1029:774], zll_main_loop72_in[1029:774], zll_main_loop72_in[773:262], zll_main_loop72_in[261:6], zll_main_loop72_in[5:0]};
  assign zll_main_loop60_in = {zll_main_loop15_in[1323:1292], zll_main_loop15_in[1291:1286], zll_main_loop15_in[1285:0]};
  assign zll_main_loop3_in = {zll_main_loop60_in[1285:1030], zll_main_loop60_in[1323:1292], zll_main_loop60_in[1291:1286], zll_main_loop60_in[1029:774], zll_main_loop60_in[773:262], zll_main_loop60_in[261:6], zll_main_loop60_in[5:0]};
  assign zll_main_loop5_in = {zll_main_loop3_in[1323:1068], zll_main_loop3_in[1067:1036], zll_main_loop3_in[773:262], zll_main_loop3_in[1035:1030], zll_main_loop3_in[1029:774], zll_main_loop3_in[261:6], zll_main_loop3_in[5:0]};
  assign zll_main_loop35_in = {zll_main_loop5_in[1067:1036], zll_main_loop5_in[523:518], zll_main_loop5_in[1323:1068], zll_main_loop5_in[517:262], zll_main_loop5_in[1035:524], zll_main_loop5_in[261:6], zll_main_loop5_in[5:0]};
  assign main_seed_in = zll_main_loop35_in[1291:1286];
  assign lit_in = main_seed_in[5:0];
  assign lit_inR1 = main_seed_in[5:0];
  assign lit_inR2 = main_seed_in[5:0];
  assign lit_inR3 = main_seed_in[5:0];
  assign lit_inR4 = main_seed_in[5:0];
  assign lit_inR5 = main_seed_in[5:0];
  assign lit_inR6 = main_seed_in[5:0];
  assign lit_inR7 = main_seed_in[5:0];
  assign lit_inR8 = main_seed_in[5:0];
  assign lit_inR9 = main_seed_in[5:0];
  assign lit_inR10 = main_seed_in[5:0];
  assign lit_inR11 = main_seed_in[5:0];
  assign lit_inR12 = main_seed_in[5:0];
  assign lit_inR13 = main_seed_in[5:0];
  assign lit_inR14 = main_seed_in[5:0];
  assign lit_inR15 = main_seed_in[5:0];
  assign lit_inR16 = main_seed_in[5:0];
  assign lit_inR17 = main_seed_in[5:0];
  assign lit_inR18 = main_seed_in[5:0];
  assign lit_inR19 = main_seed_in[5:0];
  assign lit_inR20 = main_seed_in[5:0];
  assign lit_inR21 = main_seed_in[5:0];
  assign lit_inR22 = main_seed_in[5:0];
  assign lit_inR23 = main_seed_in[5:0];
  assign lit_inR24 = main_seed_in[5:0];
  assign lit_inR25 = main_seed_in[5:0];
  assign lit_inR26 = main_seed_in[5:0];
  assign lit_inR27 = main_seed_in[5:0];
  assign lit_inR28 = main_seed_in[5:0];
  assign lit_inR29 = main_seed_in[5:0];
  assign lit_inR30 = main_seed_in[5:0];
  assign lit_inR31 = main_seed_in[5:0];
  assign lit_inR32 = main_seed_in[5:0];
  assign lit_inR33 = main_seed_in[5:0];
  assign lit_inR34 = main_seed_in[5:0];
  assign lit_inR35 = main_seed_in[5:0];
  assign lit_inR36 = main_seed_in[5:0];
  assign lit_inR37 = main_seed_in[5:0];
  assign lit_inR38 = main_seed_in[5:0];
  assign lit_inR39 = main_seed_in[5:0];
  assign lit_inR40 = main_seed_in[5:0];
  assign lit_inR41 = main_seed_in[5:0];
  assign lit_inR42 = main_seed_in[5:0];
  assign lit_inR43 = main_seed_in[5:0];
  assign lit_inR44 = main_seed_in[5:0];
  assign lit_inR45 = main_seed_in[5:0];
  assign lit_inR46 = main_seed_in[5:0];
  assign lit_inR47 = main_seed_in[5:0];
  assign lit_inR48 = main_seed_in[5:0];
  assign lit_inR49 = main_seed_in[5:0];
  assign lit_inR50 = main_seed_in[5:0];
  assign lit_inR51 = main_seed_in[5:0];
  assign lit_inR52 = main_seed_in[5:0];
  assign lit_inR53 = main_seed_in[5:0];
  assign lit_inR54 = main_seed_in[5:0];
  assign lit_inR55 = main_seed_in[5:0];
  assign lit_inR56 = main_seed_in[5:0];
  assign lit_inR57 = main_seed_in[5:0];
  assign lit_inR58 = main_seed_in[5:0];
  assign lit_inR59 = main_seed_in[5:0];
  assign lit_inR60 = main_seed_in[5:0];
  assign lit_inR61 = main_seed_in[5:0];
  assign lit_inR62 = main_seed_in[5:0];
  assign main_step256_in = {(lit_inR62[5:0] == 6'h0) ? 32'h428a2f98 : ((lit_inR61[5:0] == 6'h1) ? 32'h71374491 : ((lit_inR60[5:0] == 6'h2) ? 32'hb5c0fbcf : ((lit_inR59[5:0] == 6'h3) ? 32'he9b5dba5 : ((lit_inR58[5:0] == 6'h4) ? 32'h3956c25b : ((lit_inR57[5:0] == 6'h5) ? 32'h59f111f1 : ((lit_inR56[5:0] == 6'h6) ? 32'h923f82a4 : ((lit_inR55[5:0] == 6'h7) ? 32'hab1c5ed5 : ((lit_inR54[5:0] == 6'h8) ? 32'hd807aa98 : ((lit_inR53[5:0] == 6'h9) ? 32'h12835b01 : ((lit_inR52[5:0] == 6'ha) ? 32'h243185be : ((lit_inR51[5:0] == 6'hb) ? 32'h550c7dc3 : ((lit_inR50[5:0] == 6'hc) ? 32'h72be5d74 : ((lit_inR49[5:0] == 6'hd) ? 32'h80deb1fe : ((lit_inR48[5:0] == 6'he) ? 32'h9bdc06a7 : ((lit_inR47[5:0] == 6'hf) ? 32'hc19bf174 : ((lit_inR46[5:0] == 6'h10) ? 32'he49b69c1 : ((lit_inR45[5:0] == 6'h11) ? 32'hefbe4786 : ((lit_inR44[5:0] == 6'h12) ? 32'hfc19dc6 : ((lit_inR43[5:0] == 6'h13) ? 32'h240ca1cc : ((lit_inR42[5:0] == 6'h14) ? 32'h2de92c6f : ((lit_inR41[5:0] == 6'h15) ? 32'h4a7484aa : ((lit_inR40[5:0] == 6'h16) ? 32'h5cb0a9dc : ((lit_inR39[5:0] == 6'h17) ? 32'h76f988da : ((lit_inR38[5:0] == 6'h18) ? 32'h983e5152 : ((lit_inR37[5:0] == 6'h19) ? 32'ha831c66d : ((lit_inR36[5:0] == 6'h1a) ? 32'hb00327c8 : ((lit_inR35[5:0] == 6'h1b) ? 32'hbf597fc7 : ((lit_inR34[5:0] == 6'h1c) ? 32'hc6e00bf3 : ((lit_inR33[5:0] == 6'h1d) ? 32'hd5a79147 : ((lit_inR32[5:0] == 6'h1e) ? 32'h6ca6351 : ((lit_inR31[5:0] == 6'h1f) ? 32'h14292967 : ((lit_inR30[5:0] == 6'h20) ? 32'h27b70a85 : ((lit_inR29[5:0] == 6'h21) ? 32'h2e1b2138 : ((lit_inR28[5:0] == 6'h22) ? 32'h4d2c6dfc : ((lit_inR27[5:0] == 6'h23) ? 32'h53380d13 : ((lit_inR26[5:0] == 6'h24) ? 32'h650a7354 : ((lit_inR25[5:0] == 6'h25) ? 32'h766a0abb : ((lit_inR24[5:0] == 6'h26) ? 32'h81c2c92e : ((lit_inR23[5:0] == 6'h27) ? 32'h92722c85 : ((lit_inR22[5:0] == 6'h28) ? 32'ha2bfe8a1 : ((lit_inR21[5:0] == 6'h29) ? 32'ha81a664b : ((lit_inR20[5:0] == 6'h2a) ? 32'hc24b8b70 : ((lit_inR19[5:0] == 6'h2b) ? 32'hc76c51a3 : ((lit_inR18[5:0] == 6'h2c) ? 32'hd192e819 : ((lit_inR17[5:0] == 6'h2d) ? 32'hd6990624 : ((lit_inR16[5:0] == 6'h2e) ? 32'hf40e3585 : ((lit_inR15[5:0] == 6'h2f) ? 32'h106aa070 : ((lit_inR14[5:0] == 6'h30) ? 32'h19a4c116 : ((lit_inR13[5:0] == 6'h31) ? 32'h1e376c08 : ((lit_inR12[5:0] == 6'h32) ? 32'h2748774c : ((lit_inR11[5:0] == 6'h33) ? 32'h34b0bcb5 : ((lit_inR10[5:0] == 6'h34) ? 32'h391c0cb3 : ((lit_inR9[5:0] == 6'h35) ? 32'h4ed8aa4a : ((lit_inR8[5:0] == 6'h36) ? 32'h5b9cca4f : ((lit_inR7[5:0] == 6'h37) ? 32'h682e6ff3 : ((lit_inR6[5:0] == 6'h38) ? 32'h748f82ee : ((lit_inR5[5:0] == 6'h39) ? 32'h78a5636f : ((lit_inR4[5:0] == 6'h3a) ? 32'h84c87814 : ((lit_inR3[5:0] == 6'h3b) ? 32'h8cc70208 : ((lit_inR2[5:0] == 6'h3c) ? 32'h90befffa : ((lit_inR1[5:0] == 6'h3d) ? 32'ha4506ceb : ((lit_in[5:0] == 6'h3e) ? 32'hbef9a3f7 : 32'hc67178f2)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))), zll_main_loop35_in[1323:1292], zll_main_loop35_in[1285:1030]};
  assign zll_main_step2568_in = {main_step256_in[319:288], main_step256_in[287:256], main_step256_in[255:0]};
  assign zll_main_step2562_in = {zll_main_step2568_in[319:288], zll_main_step2568_in[255:224], zll_main_step2568_in[287:256], zll_main_step2568_in[223:192], zll_main_step2568_in[191:160], zll_main_step2568_in[159:128], zll_main_step2568_in[127:96], zll_main_step2568_in[95:64], zll_main_step2568_in[63:32], zll_main_step2568_in[31:0]};
  assign zll_main_step2561_in = {zll_main_step2562_in[319:288], zll_main_step2562_in[287:256], zll_main_step2562_in[255:224], zll_main_step2562_in[223:192], zll_main_step2562_in[159:128], zll_main_step2562_in[191:160], zll_main_step2562_in[127:96], zll_main_step2562_in[95:64], zll_main_step2562_in[63:32], zll_main_step2562_in[31:0]};
  assign zll_main_step256_in = {zll_main_step2561_in[319:288], zll_main_step2561_in[287:256], zll_main_step2561_in[255:224], zll_main_step2561_in[127:96], zll_main_step2561_in[223:192], zll_main_step2561_in[191:160], zll_main_step2561_in[159:128], zll_main_step2561_in[95:64], zll_main_step2561_in[63:32], zll_main_step2561_in[31:0]};
  assign zll_main_step2565_in = {zll_main_step256_in[319:288], zll_main_step256_in[287:256], zll_main_step256_in[255:224], zll_main_step256_in[223:192], zll_main_step256_in[191:160], zll_main_step256_in[159:128], zll_main_step256_in[95:64], zll_main_step256_in[127:96], zll_main_step256_in[63:32], zll_main_step256_in[31:0]};
  assign zll_main_step2566_in = {zll_main_step2565_in[319:288], zll_main_step2565_in[287:256], zll_main_step2565_in[255:224], zll_main_step2565_in[63:32], zll_main_step2565_in[223:192], zll_main_step2565_in[191:160], zll_main_step2565_in[159:128], zll_main_step2565_in[127:96], zll_main_step2565_in[95:64], zll_main_step2565_in[31:0]};
  assign main_bigsigma1_in = zll_main_step2566_in[191:160];
  Main_bigsigma1  instR7 (main_bigsigma1_in[31:0], main_bigsigma1_out);
  assign main_ch_in = {zll_main_step2566_in[191:160], zll_main_step2566_in[95:64], zll_main_step2566_in[223:192]};
  Main_ch  instR8 (main_ch_in[95:64], main_ch_in[63:32], main_ch_in[31:0], main_ch_out);
  assign plusw32_inR3 = {main_bigsigma1_out, main_ch_out};
  plusW32  instR9 (plusw32_inR3[63:32], plusw32_inR3[31:0], extresR7[31:0]);
  assign plusw32_inR4 = {zll_main_step2566_in[319:288], zll_main_step2566_in[255:224]};
  plusW32  instR10 (plusw32_inR4[63:32], plusw32_inR4[31:0], extresR8[31:0]);
  assign plusw32_inR5 = {extresR7, extresR8};
  plusW32  instR11 (plusw32_inR5[63:32], plusw32_inR5[31:0], extresR9[31:0]);
  assign plusw32_inR6 = {zll_main_step2566_in[31:0], extresR9};
  plusW32  instR12 (plusw32_inR6[63:32], plusw32_inR6[31:0], extresR10[31:0]);
  assign main_bigsigma0_in = zll_main_step2566_in[287:256];
  assign main_rotater2_in = main_bigsigma0_in[31:0];
  assign zll_main_rotater211_in = main_rotater2_in[31:0];
  assign zll_main_rotater210_in = {zll_main_rotater211_in[30], zll_main_rotater211_in[31], zll_main_rotater211_in[29], zll_main_rotater211_in[28], zll_main_rotater211_in[27], zll_main_rotater211_in[26], zll_main_rotater211_in[25], zll_main_rotater211_in[24], zll_main_rotater211_in[23], zll_main_rotater211_in[22], zll_main_rotater211_in[21], zll_main_rotater211_in[20], zll_main_rotater211_in[19], zll_main_rotater211_in[18], zll_main_rotater211_in[17], zll_main_rotater211_in[16], zll_main_rotater211_in[15], zll_main_rotater211_in[14], zll_main_rotater211_in[13], zll_main_rotater211_in[12], zll_main_rotater211_in[11], zll_main_rotater211_in[10], zll_main_rotater211_in[9], zll_main_rotater211_in[8], zll_main_rotater211_in[7], zll_main_rotater211_in[6], zll_main_rotater211_in[5], zll_main_rotater211_in[4], zll_main_rotater211_in[3], zll_main_rotater211_in[2], zll_main_rotater211_in[1], zll_main_rotater211_in[0]};
  assign zll_main_rotater213_in = {zll_main_rotater210_in[31], zll_main_rotater210_in[29], zll_main_rotater210_in[30], zll_main_rotater210_in[28], zll_main_rotater210_in[27], zll_main_rotater210_in[26], zll_main_rotater210_in[25], zll_main_rotater210_in[24], zll_main_rotater210_in[23], zll_main_rotater210_in[22], zll_main_rotater210_in[21], zll_main_rotater210_in[20], zll_main_rotater210_in[19], zll_main_rotater210_in[18], zll_main_rotater210_in[17], zll_main_rotater210_in[16], zll_main_rotater210_in[15], zll_main_rotater210_in[14], zll_main_rotater210_in[13], zll_main_rotater210_in[12], zll_main_rotater210_in[11], zll_main_rotater210_in[10], zll_main_rotater210_in[9], zll_main_rotater210_in[8], zll_main_rotater210_in[7], zll_main_rotater210_in[6], zll_main_rotater210_in[5], zll_main_rotater210_in[4], zll_main_rotater210_in[3], zll_main_rotater210_in[2], zll_main_rotater210_in[1], zll_main_rotater210_in[0]};
  assign zll_main_rotater23_in = {zll_main_rotater213_in[31], zll_main_rotater213_in[27], zll_main_rotater213_in[30], zll_main_rotater213_in[29], zll_main_rotater213_in[28], zll_main_rotater213_in[26], zll_main_rotater213_in[25], zll_main_rotater213_in[24], zll_main_rotater213_in[23], zll_main_rotater213_in[22], zll_main_rotater213_in[21], zll_main_rotater213_in[20], zll_main_rotater213_in[19], zll_main_rotater213_in[18], zll_main_rotater213_in[17], zll_main_rotater213_in[16], zll_main_rotater213_in[15], zll_main_rotater213_in[14], zll_main_rotater213_in[13], zll_main_rotater213_in[12], zll_main_rotater213_in[11], zll_main_rotater213_in[10], zll_main_rotater213_in[9], zll_main_rotater213_in[8], zll_main_rotater213_in[7], zll_main_rotater213_in[6], zll_main_rotater213_in[5], zll_main_rotater213_in[4], zll_main_rotater213_in[3], zll_main_rotater213_in[2], zll_main_rotater213_in[1], zll_main_rotater213_in[0]};
  assign zll_main_rotater242_in = {zll_main_rotater23_in[26], zll_main_rotater23_in[31], zll_main_rotater23_in[30], zll_main_rotater23_in[29], zll_main_rotater23_in[28], zll_main_rotater23_in[27], zll_main_rotater23_in[25], zll_main_rotater23_in[24], zll_main_rotater23_in[23], zll_main_rotater23_in[22], zll_main_rotater23_in[21], zll_main_rotater23_in[20], zll_main_rotater23_in[19], zll_main_rotater23_in[18], zll_main_rotater23_in[17], zll_main_rotater23_in[16], zll_main_rotater23_in[15], zll_main_rotater23_in[14], zll_main_rotater23_in[13], zll_main_rotater23_in[12], zll_main_rotater23_in[11], zll_main_rotater23_in[10], zll_main_rotater23_in[9], zll_main_rotater23_in[8], zll_main_rotater23_in[7], zll_main_rotater23_in[6], zll_main_rotater23_in[5], zll_main_rotater23_in[4], zll_main_rotater23_in[3], zll_main_rotater23_in[2], zll_main_rotater23_in[1], zll_main_rotater23_in[0]};
  assign zll_main_rotater220_in = {zll_main_rotater242_in[31], zll_main_rotater242_in[25], zll_main_rotater242_in[30], zll_main_rotater242_in[29], zll_main_rotater242_in[28], zll_main_rotater242_in[27], zll_main_rotater242_in[26], zll_main_rotater242_in[24], zll_main_rotater242_in[23], zll_main_rotater242_in[22], zll_main_rotater242_in[21], zll_main_rotater242_in[20], zll_main_rotater242_in[19], zll_main_rotater242_in[18], zll_main_rotater242_in[17], zll_main_rotater242_in[16], zll_main_rotater242_in[15], zll_main_rotater242_in[14], zll_main_rotater242_in[13], zll_main_rotater242_in[12], zll_main_rotater242_in[11], zll_main_rotater242_in[10], zll_main_rotater242_in[9], zll_main_rotater242_in[8], zll_main_rotater242_in[7], zll_main_rotater242_in[6], zll_main_rotater242_in[5], zll_main_rotater242_in[4], zll_main_rotater242_in[3], zll_main_rotater242_in[2], zll_main_rotater242_in[1], zll_main_rotater242_in[0]};
  assign zll_main_rotater24_in = {zll_main_rotater220_in[31], zll_main_rotater220_in[30], zll_main_rotater220_in[29], zll_main_rotater220_in[28], zll_main_rotater220_in[27], zll_main_rotater220_in[24], zll_main_rotater220_in[26], zll_main_rotater220_in[25], zll_main_rotater220_in[23], zll_main_rotater220_in[22], zll_main_rotater220_in[21], zll_main_rotater220_in[20], zll_main_rotater220_in[19], zll_main_rotater220_in[18], zll_main_rotater220_in[17], zll_main_rotater220_in[16], zll_main_rotater220_in[15], zll_main_rotater220_in[14], zll_main_rotater220_in[13], zll_main_rotater220_in[12], zll_main_rotater220_in[11], zll_main_rotater220_in[10], zll_main_rotater220_in[9], zll_main_rotater220_in[8], zll_main_rotater220_in[7], zll_main_rotater220_in[6], zll_main_rotater220_in[5], zll_main_rotater220_in[4], zll_main_rotater220_in[3], zll_main_rotater220_in[2], zll_main_rotater220_in[1], zll_main_rotater220_in[0]};
  assign zll_main_rotater233_in = {zll_main_rotater24_in[31], zll_main_rotater24_in[30], zll_main_rotater24_in[29], zll_main_rotater24_in[28], zll_main_rotater24_in[23], zll_main_rotater24_in[27], zll_main_rotater24_in[26], zll_main_rotater24_in[25], zll_main_rotater24_in[24], zll_main_rotater24_in[22], zll_main_rotater24_in[21], zll_main_rotater24_in[20], zll_main_rotater24_in[19], zll_main_rotater24_in[18], zll_main_rotater24_in[17], zll_main_rotater24_in[16], zll_main_rotater24_in[15], zll_main_rotater24_in[14], zll_main_rotater24_in[13], zll_main_rotater24_in[12], zll_main_rotater24_in[11], zll_main_rotater24_in[10], zll_main_rotater24_in[9], zll_main_rotater24_in[8], zll_main_rotater24_in[7], zll_main_rotater24_in[6], zll_main_rotater24_in[5], zll_main_rotater24_in[4], zll_main_rotater24_in[3], zll_main_rotater24_in[2], zll_main_rotater24_in[1], zll_main_rotater24_in[0]};
  assign zll_main_rotater212_in = {zll_main_rotater233_in[31], zll_main_rotater233_in[30], zll_main_rotater233_in[29], zll_main_rotater233_in[28], zll_main_rotater233_in[27], zll_main_rotater233_in[22], zll_main_rotater233_in[26], zll_main_rotater233_in[25], zll_main_rotater233_in[24], zll_main_rotater233_in[23], zll_main_rotater233_in[21], zll_main_rotater233_in[20], zll_main_rotater233_in[19], zll_main_rotater233_in[18], zll_main_rotater233_in[17], zll_main_rotater233_in[16], zll_main_rotater233_in[15], zll_main_rotater233_in[14], zll_main_rotater233_in[13], zll_main_rotater233_in[12], zll_main_rotater233_in[11], zll_main_rotater233_in[10], zll_main_rotater233_in[9], zll_main_rotater233_in[8], zll_main_rotater233_in[7], zll_main_rotater233_in[6], zll_main_rotater233_in[5], zll_main_rotater233_in[4], zll_main_rotater233_in[3], zll_main_rotater233_in[2], zll_main_rotater233_in[1], zll_main_rotater233_in[0]};
  assign zll_main_rotater235_in = {zll_main_rotater212_in[21], zll_main_rotater212_in[31], zll_main_rotater212_in[30], zll_main_rotater212_in[29], zll_main_rotater212_in[28], zll_main_rotater212_in[27], zll_main_rotater212_in[26], zll_main_rotater212_in[25], zll_main_rotater212_in[24], zll_main_rotater212_in[23], zll_main_rotater212_in[22], zll_main_rotater212_in[20], zll_main_rotater212_in[19], zll_main_rotater212_in[18], zll_main_rotater212_in[17], zll_main_rotater212_in[16], zll_main_rotater212_in[15], zll_main_rotater212_in[14], zll_main_rotater212_in[13], zll_main_rotater212_in[12], zll_main_rotater212_in[11], zll_main_rotater212_in[10], zll_main_rotater212_in[9], zll_main_rotater212_in[8], zll_main_rotater212_in[7], zll_main_rotater212_in[6], zll_main_rotater212_in[5], zll_main_rotater212_in[4], zll_main_rotater212_in[3], zll_main_rotater212_in[2], zll_main_rotater212_in[1], zll_main_rotater212_in[0]};
  assign zll_main_rotater230_in = {zll_main_rotater235_in[31], zll_main_rotater235_in[30], zll_main_rotater235_in[20], zll_main_rotater235_in[29], zll_main_rotater235_in[28], zll_main_rotater235_in[27], zll_main_rotater235_in[26], zll_main_rotater235_in[25], zll_main_rotater235_in[24], zll_main_rotater235_in[23], zll_main_rotater235_in[22], zll_main_rotater235_in[21], zll_main_rotater235_in[19], zll_main_rotater235_in[18], zll_main_rotater235_in[17], zll_main_rotater235_in[16], zll_main_rotater235_in[15], zll_main_rotater235_in[14], zll_main_rotater235_in[13], zll_main_rotater235_in[12], zll_main_rotater235_in[11], zll_main_rotater235_in[10], zll_main_rotater235_in[9], zll_main_rotater235_in[8], zll_main_rotater235_in[7], zll_main_rotater235_in[6], zll_main_rotater235_in[5], zll_main_rotater235_in[4], zll_main_rotater235_in[3], zll_main_rotater235_in[2], zll_main_rotater235_in[1], zll_main_rotater235_in[0]};
  assign zll_main_rotater26_in = {zll_main_rotater230_in[31], zll_main_rotater230_in[30], zll_main_rotater230_in[29], zll_main_rotater230_in[28], zll_main_rotater230_in[27], zll_main_rotater230_in[26], zll_main_rotater230_in[19], zll_main_rotater230_in[25], zll_main_rotater230_in[24], zll_main_rotater230_in[23], zll_main_rotater230_in[22], zll_main_rotater230_in[21], zll_main_rotater230_in[20], zll_main_rotater230_in[18], zll_main_rotater230_in[17], zll_main_rotater230_in[16], zll_main_rotater230_in[15], zll_main_rotater230_in[14], zll_main_rotater230_in[13], zll_main_rotater230_in[12], zll_main_rotater230_in[11], zll_main_rotater230_in[10], zll_main_rotater230_in[9], zll_main_rotater230_in[8], zll_main_rotater230_in[7], zll_main_rotater230_in[6], zll_main_rotater230_in[5], zll_main_rotater230_in[4], zll_main_rotater230_in[3], zll_main_rotater230_in[2], zll_main_rotater230_in[1], zll_main_rotater230_in[0]};
  assign zll_main_rotater232_in = {zll_main_rotater26_in[31], zll_main_rotater26_in[18], zll_main_rotater26_in[30], zll_main_rotater26_in[29], zll_main_rotater26_in[28], zll_main_rotater26_in[27], zll_main_rotater26_in[26], zll_main_rotater26_in[25], zll_main_rotater26_in[24], zll_main_rotater26_in[23], zll_main_rotater26_in[22], zll_main_rotater26_in[21], zll_main_rotater26_in[20], zll_main_rotater26_in[19], zll_main_rotater26_in[17], zll_main_rotater26_in[16], zll_main_rotater26_in[15], zll_main_rotater26_in[14], zll_main_rotater26_in[13], zll_main_rotater26_in[12], zll_main_rotater26_in[11], zll_main_rotater26_in[10], zll_main_rotater26_in[9], zll_main_rotater26_in[8], zll_main_rotater26_in[7], zll_main_rotater26_in[6], zll_main_rotater26_in[5], zll_main_rotater26_in[4], zll_main_rotater26_in[3], zll_main_rotater26_in[2], zll_main_rotater26_in[1], zll_main_rotater26_in[0]};
  assign zll_main_rotater236_in = {zll_main_rotater232_in[31], zll_main_rotater232_in[30], zll_main_rotater232_in[29], zll_main_rotater232_in[28], zll_main_rotater232_in[17], zll_main_rotater232_in[27], zll_main_rotater232_in[26], zll_main_rotater232_in[25], zll_main_rotater232_in[24], zll_main_rotater232_in[23], zll_main_rotater232_in[22], zll_main_rotater232_in[21], zll_main_rotater232_in[20], zll_main_rotater232_in[19], zll_main_rotater232_in[18], zll_main_rotater232_in[16], zll_main_rotater232_in[15], zll_main_rotater232_in[14], zll_main_rotater232_in[13], zll_main_rotater232_in[12], zll_main_rotater232_in[11], zll_main_rotater232_in[10], zll_main_rotater232_in[9], zll_main_rotater232_in[8], zll_main_rotater232_in[7], zll_main_rotater232_in[6], zll_main_rotater232_in[5], zll_main_rotater232_in[4], zll_main_rotater232_in[3], zll_main_rotater232_in[2], zll_main_rotater232_in[1], zll_main_rotater232_in[0]};
  assign zll_main_rotater216_in = {zll_main_rotater236_in[31], zll_main_rotater236_in[30], zll_main_rotater236_in[29], zll_main_rotater236_in[28], zll_main_rotater236_in[27], zll_main_rotater236_in[26], zll_main_rotater236_in[25], zll_main_rotater236_in[24], zll_main_rotater236_in[23], zll_main_rotater236_in[22], zll_main_rotater236_in[21], zll_main_rotater236_in[20], zll_main_rotater236_in[19], zll_main_rotater236_in[16], zll_main_rotater236_in[18], zll_main_rotater236_in[17], zll_main_rotater236_in[15], zll_main_rotater236_in[14], zll_main_rotater236_in[13], zll_main_rotater236_in[12], zll_main_rotater236_in[11], zll_main_rotater236_in[10], zll_main_rotater236_in[9], zll_main_rotater236_in[8], zll_main_rotater236_in[7], zll_main_rotater236_in[6], zll_main_rotater236_in[5], zll_main_rotater236_in[4], zll_main_rotater236_in[3], zll_main_rotater236_in[2], zll_main_rotater236_in[1], zll_main_rotater236_in[0]};
  assign zll_main_rotater241_in = {zll_main_rotater216_in[31], zll_main_rotater216_in[30], zll_main_rotater216_in[29], zll_main_rotater216_in[15], zll_main_rotater216_in[28], zll_main_rotater216_in[27], zll_main_rotater216_in[26], zll_main_rotater216_in[25], zll_main_rotater216_in[24], zll_main_rotater216_in[23], zll_main_rotater216_in[22], zll_main_rotater216_in[21], zll_main_rotater216_in[20], zll_main_rotater216_in[19], zll_main_rotater216_in[18], zll_main_rotater216_in[17], zll_main_rotater216_in[16], zll_main_rotater216_in[14], zll_main_rotater216_in[13], zll_main_rotater216_in[12], zll_main_rotater216_in[11], zll_main_rotater216_in[10], zll_main_rotater216_in[9], zll_main_rotater216_in[8], zll_main_rotater216_in[7], zll_main_rotater216_in[6], zll_main_rotater216_in[5], zll_main_rotater216_in[4], zll_main_rotater216_in[3], zll_main_rotater216_in[2], zll_main_rotater216_in[1], zll_main_rotater216_in[0]};
  assign zll_main_rotater29_in = {zll_main_rotater241_in[31], zll_main_rotater241_in[30], zll_main_rotater241_in[29], zll_main_rotater241_in[28], zll_main_rotater241_in[27], zll_main_rotater241_in[26], zll_main_rotater241_in[25], zll_main_rotater241_in[14], zll_main_rotater241_in[24], zll_main_rotater241_in[23], zll_main_rotater241_in[22], zll_main_rotater241_in[21], zll_main_rotater241_in[20], zll_main_rotater241_in[19], zll_main_rotater241_in[18], zll_main_rotater241_in[17], zll_main_rotater241_in[16], zll_main_rotater241_in[15], zll_main_rotater241_in[13], zll_main_rotater241_in[12], zll_main_rotater241_in[11], zll_main_rotater241_in[10], zll_main_rotater241_in[9], zll_main_rotater241_in[8], zll_main_rotater241_in[7], zll_main_rotater241_in[6], zll_main_rotater241_in[5], zll_main_rotater241_in[4], zll_main_rotater241_in[3], zll_main_rotater241_in[2], zll_main_rotater241_in[1], zll_main_rotater241_in[0]};
  assign zll_main_rotater218_in = {zll_main_rotater29_in[31], zll_main_rotater29_in[30], zll_main_rotater29_in[29], zll_main_rotater29_in[28], zll_main_rotater29_in[27], zll_main_rotater29_in[26], zll_main_rotater29_in[25], zll_main_rotater29_in[24], zll_main_rotater29_in[12], zll_main_rotater29_in[23], zll_main_rotater29_in[22], zll_main_rotater29_in[21], zll_main_rotater29_in[20], zll_main_rotater29_in[19], zll_main_rotater29_in[18], zll_main_rotater29_in[17], zll_main_rotater29_in[16], zll_main_rotater29_in[15], zll_main_rotater29_in[14], zll_main_rotater29_in[13], zll_main_rotater29_in[11], zll_main_rotater29_in[10], zll_main_rotater29_in[9], zll_main_rotater29_in[8], zll_main_rotater29_in[7], zll_main_rotater29_in[6], zll_main_rotater29_in[5], zll_main_rotater29_in[4], zll_main_rotater29_in[3], zll_main_rotater29_in[2], zll_main_rotater29_in[1], zll_main_rotater29_in[0]};
  assign zll_main_rotater239_in = {zll_main_rotater218_in[31], zll_main_rotater218_in[30], zll_main_rotater218_in[29], zll_main_rotater218_in[28], zll_main_rotater218_in[27], zll_main_rotater218_in[26], zll_main_rotater218_in[25], zll_main_rotater218_in[24], zll_main_rotater218_in[23], zll_main_rotater218_in[22], zll_main_rotater218_in[21], zll_main_rotater218_in[20], zll_main_rotater218_in[19], zll_main_rotater218_in[18], zll_main_rotater218_in[17], zll_main_rotater218_in[16], zll_main_rotater218_in[15], zll_main_rotater218_in[14], zll_main_rotater218_in[11], zll_main_rotater218_in[13], zll_main_rotater218_in[12], zll_main_rotater218_in[10], zll_main_rotater218_in[9], zll_main_rotater218_in[8], zll_main_rotater218_in[7], zll_main_rotater218_in[6], zll_main_rotater218_in[5], zll_main_rotater218_in[4], zll_main_rotater218_in[3], zll_main_rotater218_in[2], zll_main_rotater218_in[1], zll_main_rotater218_in[0]};
  assign zll_main_rotater231_in = {zll_main_rotater239_in[31], zll_main_rotater239_in[30], zll_main_rotater239_in[29], zll_main_rotater239_in[28], zll_main_rotater239_in[27], zll_main_rotater239_in[26], zll_main_rotater239_in[25], zll_main_rotater239_in[24], zll_main_rotater239_in[23], zll_main_rotater239_in[22], zll_main_rotater239_in[21], zll_main_rotater239_in[20], zll_main_rotater239_in[19], zll_main_rotater239_in[18], zll_main_rotater239_in[10], zll_main_rotater239_in[17], zll_main_rotater239_in[16], zll_main_rotater239_in[15], zll_main_rotater239_in[14], zll_main_rotater239_in[13], zll_main_rotater239_in[12], zll_main_rotater239_in[11], zll_main_rotater239_in[9], zll_main_rotater239_in[8], zll_main_rotater239_in[7], zll_main_rotater239_in[6], zll_main_rotater239_in[5], zll_main_rotater239_in[4], zll_main_rotater239_in[3], zll_main_rotater239_in[2], zll_main_rotater239_in[1], zll_main_rotater239_in[0]};
  assign zll_main_rotater28_in = {zll_main_rotater231_in[31], zll_main_rotater231_in[30], zll_main_rotater231_in[29], zll_main_rotater231_in[28], zll_main_rotater231_in[27], zll_main_rotater231_in[26], zll_main_rotater231_in[25], zll_main_rotater231_in[24], zll_main_rotater231_in[23], zll_main_rotater231_in[22], zll_main_rotater231_in[21], zll_main_rotater231_in[20], zll_main_rotater231_in[19], zll_main_rotater231_in[18], zll_main_rotater231_in[17], zll_main_rotater231_in[16], zll_main_rotater231_in[15], zll_main_rotater231_in[14], zll_main_rotater231_in[13], zll_main_rotater231_in[9], zll_main_rotater231_in[12], zll_main_rotater231_in[11], zll_main_rotater231_in[10], zll_main_rotater231_in[8], zll_main_rotater231_in[7], zll_main_rotater231_in[6], zll_main_rotater231_in[5], zll_main_rotater231_in[4], zll_main_rotater231_in[3], zll_main_rotater231_in[2], zll_main_rotater231_in[1], zll_main_rotater231_in[0]};
  assign zll_main_rotater215_in = {zll_main_rotater28_in[31], zll_main_rotater28_in[30], zll_main_rotater28_in[29], zll_main_rotater28_in[28], zll_main_rotater28_in[27], zll_main_rotater28_in[26], zll_main_rotater28_in[25], zll_main_rotater28_in[24], zll_main_rotater28_in[23], zll_main_rotater28_in[22], zll_main_rotater28_in[21], zll_main_rotater28_in[20], zll_main_rotater28_in[19], zll_main_rotater28_in[18], zll_main_rotater28_in[17], zll_main_rotater28_in[16], zll_main_rotater28_in[15], zll_main_rotater28_in[14], zll_main_rotater28_in[13], zll_main_rotater28_in[8], zll_main_rotater28_in[12], zll_main_rotater28_in[11], zll_main_rotater28_in[10], zll_main_rotater28_in[9], zll_main_rotater28_in[7], zll_main_rotater28_in[6], zll_main_rotater28_in[5], zll_main_rotater28_in[4], zll_main_rotater28_in[3], zll_main_rotater28_in[2], zll_main_rotater28_in[1], zll_main_rotater28_in[0]};
  assign zll_main_rotater219_in = {zll_main_rotater215_in[31], zll_main_rotater215_in[30], zll_main_rotater215_in[29], zll_main_rotater215_in[28], zll_main_rotater215_in[27], zll_main_rotater215_in[26], zll_main_rotater215_in[25], zll_main_rotater215_in[24], zll_main_rotater215_in[7], zll_main_rotater215_in[23], zll_main_rotater215_in[22], zll_main_rotater215_in[21], zll_main_rotater215_in[20], zll_main_rotater215_in[19], zll_main_rotater215_in[18], zll_main_rotater215_in[17], zll_main_rotater215_in[16], zll_main_rotater215_in[15], zll_main_rotater215_in[14], zll_main_rotater215_in[13], zll_main_rotater215_in[12], zll_main_rotater215_in[11], zll_main_rotater215_in[10], zll_main_rotater215_in[9], zll_main_rotater215_in[8], zll_main_rotater215_in[6], zll_main_rotater215_in[5], zll_main_rotater215_in[4], zll_main_rotater215_in[3], zll_main_rotater215_in[2], zll_main_rotater215_in[1], zll_main_rotater215_in[0]};
  assign zll_main_rotater27_in = {zll_main_rotater219_in[31], zll_main_rotater219_in[6], zll_main_rotater219_in[30], zll_main_rotater219_in[29], zll_main_rotater219_in[28], zll_main_rotater219_in[27], zll_main_rotater219_in[26], zll_main_rotater219_in[25], zll_main_rotater219_in[24], zll_main_rotater219_in[23], zll_main_rotater219_in[22], zll_main_rotater219_in[21], zll_main_rotater219_in[20], zll_main_rotater219_in[19], zll_main_rotater219_in[18], zll_main_rotater219_in[17], zll_main_rotater219_in[16], zll_main_rotater219_in[15], zll_main_rotater219_in[14], zll_main_rotater219_in[13], zll_main_rotater219_in[12], zll_main_rotater219_in[11], zll_main_rotater219_in[10], zll_main_rotater219_in[9], zll_main_rotater219_in[8], zll_main_rotater219_in[7], zll_main_rotater219_in[5], zll_main_rotater219_in[4], zll_main_rotater219_in[3], zll_main_rotater219_in[2], zll_main_rotater219_in[1], zll_main_rotater219_in[0]};
  assign zll_main_rotater214_in = {zll_main_rotater27_in[31], zll_main_rotater27_in[30], zll_main_rotater27_in[29], zll_main_rotater27_in[28], zll_main_rotater27_in[27], zll_main_rotater27_in[26], zll_main_rotater27_in[25], zll_main_rotater27_in[5], zll_main_rotater27_in[24], zll_main_rotater27_in[23], zll_main_rotater27_in[22], zll_main_rotater27_in[21], zll_main_rotater27_in[20], zll_main_rotater27_in[19], zll_main_rotater27_in[18], zll_main_rotater27_in[17], zll_main_rotater27_in[16], zll_main_rotater27_in[15], zll_main_rotater27_in[14], zll_main_rotater27_in[13], zll_main_rotater27_in[12], zll_main_rotater27_in[11], zll_main_rotater27_in[10], zll_main_rotater27_in[9], zll_main_rotater27_in[8], zll_main_rotater27_in[7], zll_main_rotater27_in[6], zll_main_rotater27_in[4], zll_main_rotater27_in[3], zll_main_rotater27_in[2], zll_main_rotater27_in[1], zll_main_rotater27_in[0]};
  assign zll_main_rotater217_in = {zll_main_rotater214_in[31], zll_main_rotater214_in[30], zll_main_rotater214_in[29], zll_main_rotater214_in[28], zll_main_rotater214_in[27], zll_main_rotater214_in[26], zll_main_rotater214_in[25], zll_main_rotater214_in[24], zll_main_rotater214_in[23], zll_main_rotater214_in[22], zll_main_rotater214_in[21], zll_main_rotater214_in[20], zll_main_rotater214_in[19], zll_main_rotater214_in[18], zll_main_rotater214_in[17], zll_main_rotater214_in[16], zll_main_rotater214_in[15], zll_main_rotater214_in[14], zll_main_rotater214_in[13], zll_main_rotater214_in[12], zll_main_rotater214_in[11], zll_main_rotater214_in[10], zll_main_rotater214_in[9], zll_main_rotater214_in[8], zll_main_rotater214_in[7], zll_main_rotater214_in[6], zll_main_rotater214_in[4], zll_main_rotater214_in[5], zll_main_rotater214_in[3], zll_main_rotater214_in[2], zll_main_rotater214_in[1], zll_main_rotater214_in[0]};
  assign zll_main_rotater240_in = {zll_main_rotater217_in[31], zll_main_rotater217_in[30], zll_main_rotater217_in[29], zll_main_rotater217_in[28], zll_main_rotater217_in[27], zll_main_rotater217_in[26], zll_main_rotater217_in[25], zll_main_rotater217_in[24], zll_main_rotater217_in[23], zll_main_rotater217_in[22], zll_main_rotater217_in[21], zll_main_rotater217_in[20], zll_main_rotater217_in[19], zll_main_rotater217_in[18], zll_main_rotater217_in[17], zll_main_rotater217_in[16], zll_main_rotater217_in[15], zll_main_rotater217_in[14], zll_main_rotater217_in[13], zll_main_rotater217_in[12], zll_main_rotater217_in[11], zll_main_rotater217_in[10], zll_main_rotater217_in[3], zll_main_rotater217_in[9], zll_main_rotater217_in[8], zll_main_rotater217_in[7], zll_main_rotater217_in[6], zll_main_rotater217_in[5], zll_main_rotater217_in[4], zll_main_rotater217_in[2], zll_main_rotater217_in[1], zll_main_rotater217_in[0]};
  assign zll_main_rotater2_in = {zll_main_rotater240_in[31], zll_main_rotater240_in[30], zll_main_rotater240_in[29], zll_main_rotater240_in[28], zll_main_rotater240_in[27], zll_main_rotater240_in[26], zll_main_rotater240_in[25], zll_main_rotater240_in[24], zll_main_rotater240_in[23], zll_main_rotater240_in[22], zll_main_rotater240_in[21], zll_main_rotater240_in[20], zll_main_rotater240_in[19], zll_main_rotater240_in[18], zll_main_rotater240_in[17], zll_main_rotater240_in[2], zll_main_rotater240_in[16], zll_main_rotater240_in[15], zll_main_rotater240_in[14], zll_main_rotater240_in[13], zll_main_rotater240_in[12], zll_main_rotater240_in[11], zll_main_rotater240_in[10], zll_main_rotater240_in[9], zll_main_rotater240_in[8], zll_main_rotater240_in[7], zll_main_rotater240_in[6], zll_main_rotater240_in[5], zll_main_rotater240_in[4], zll_main_rotater240_in[3], zll_main_rotater240_in[1], zll_main_rotater240_in[0]};
  assign zll_main_rotater237_in = {zll_main_rotater2_in[31], zll_main_rotater2_in[30], zll_main_rotater2_in[29], zll_main_rotater2_in[28], zll_main_rotater2_in[1], zll_main_rotater2_in[27], zll_main_rotater2_in[26], zll_main_rotater2_in[25], zll_main_rotater2_in[24], zll_main_rotater2_in[23], zll_main_rotater2_in[22], zll_main_rotater2_in[21], zll_main_rotater2_in[20], zll_main_rotater2_in[19], zll_main_rotater2_in[18], zll_main_rotater2_in[17], zll_main_rotater2_in[16], zll_main_rotater2_in[15], zll_main_rotater2_in[14], zll_main_rotater2_in[13], zll_main_rotater2_in[12], zll_main_rotater2_in[11], zll_main_rotater2_in[10], zll_main_rotater2_in[9], zll_main_rotater2_in[8], zll_main_rotater2_in[7], zll_main_rotater2_in[6], zll_main_rotater2_in[5], zll_main_rotater2_in[4], zll_main_rotater2_in[3], zll_main_rotater2_in[2], zll_main_rotater2_in[0]};
  assign main_rotater13_in = main_bigsigma0_in[31:0];
  assign zll_main_rotater1323_in = main_rotater13_in[31:0];
  assign zll_main_rotater1316_in = {zll_main_rotater1323_in[29], zll_main_rotater1323_in[31], zll_main_rotater1323_in[30], zll_main_rotater1323_in[28], zll_main_rotater1323_in[27], zll_main_rotater1323_in[26], zll_main_rotater1323_in[25], zll_main_rotater1323_in[24], zll_main_rotater1323_in[23], zll_main_rotater1323_in[22], zll_main_rotater1323_in[21], zll_main_rotater1323_in[20], zll_main_rotater1323_in[19], zll_main_rotater1323_in[18], zll_main_rotater1323_in[17], zll_main_rotater1323_in[16], zll_main_rotater1323_in[15], zll_main_rotater1323_in[14], zll_main_rotater1323_in[13], zll_main_rotater1323_in[12], zll_main_rotater1323_in[11], zll_main_rotater1323_in[10], zll_main_rotater1323_in[9], zll_main_rotater1323_in[8], zll_main_rotater1323_in[7], zll_main_rotater1323_in[6], zll_main_rotater1323_in[5], zll_main_rotater1323_in[4], zll_main_rotater1323_in[3], zll_main_rotater1323_in[2], zll_main_rotater1323_in[1], zll_main_rotater1323_in[0]};
  assign zll_main_rotater1328_in = {zll_main_rotater1316_in[31], zll_main_rotater1316_in[30], zll_main_rotater1316_in[28], zll_main_rotater1316_in[29], zll_main_rotater1316_in[27], zll_main_rotater1316_in[26], zll_main_rotater1316_in[25], zll_main_rotater1316_in[24], zll_main_rotater1316_in[23], zll_main_rotater1316_in[22], zll_main_rotater1316_in[21], zll_main_rotater1316_in[20], zll_main_rotater1316_in[19], zll_main_rotater1316_in[18], zll_main_rotater1316_in[17], zll_main_rotater1316_in[16], zll_main_rotater1316_in[15], zll_main_rotater1316_in[14], zll_main_rotater1316_in[13], zll_main_rotater1316_in[12], zll_main_rotater1316_in[11], zll_main_rotater1316_in[10], zll_main_rotater1316_in[9], zll_main_rotater1316_in[8], zll_main_rotater1316_in[7], zll_main_rotater1316_in[6], zll_main_rotater1316_in[5], zll_main_rotater1316_in[4], zll_main_rotater1316_in[3], zll_main_rotater1316_in[2], zll_main_rotater1316_in[1], zll_main_rotater1316_in[0]};
  assign zll_main_rotater1317_in = {zll_main_rotater1328_in[31], zll_main_rotater1328_in[30], zll_main_rotater1328_in[29], zll_main_rotater1328_in[27], zll_main_rotater1328_in[28], zll_main_rotater1328_in[26], zll_main_rotater1328_in[25], zll_main_rotater1328_in[24], zll_main_rotater1328_in[23], zll_main_rotater1328_in[22], zll_main_rotater1328_in[21], zll_main_rotater1328_in[20], zll_main_rotater1328_in[19], zll_main_rotater1328_in[18], zll_main_rotater1328_in[17], zll_main_rotater1328_in[16], zll_main_rotater1328_in[15], zll_main_rotater1328_in[14], zll_main_rotater1328_in[13], zll_main_rotater1328_in[12], zll_main_rotater1328_in[11], zll_main_rotater1328_in[10], zll_main_rotater1328_in[9], zll_main_rotater1328_in[8], zll_main_rotater1328_in[7], zll_main_rotater1328_in[6], zll_main_rotater1328_in[5], zll_main_rotater1328_in[4], zll_main_rotater1328_in[3], zll_main_rotater1328_in[2], zll_main_rotater1328_in[1], zll_main_rotater1328_in[0]};
  assign zll_main_rotater1321_in = {zll_main_rotater1317_in[31], zll_main_rotater1317_in[30], zll_main_rotater1317_in[29], zll_main_rotater1317_in[28], zll_main_rotater1317_in[26], zll_main_rotater1317_in[27], zll_main_rotater1317_in[25], zll_main_rotater1317_in[24], zll_main_rotater1317_in[23], zll_main_rotater1317_in[22], zll_main_rotater1317_in[21], zll_main_rotater1317_in[20], zll_main_rotater1317_in[19], zll_main_rotater1317_in[18], zll_main_rotater1317_in[17], zll_main_rotater1317_in[16], zll_main_rotater1317_in[15], zll_main_rotater1317_in[14], zll_main_rotater1317_in[13], zll_main_rotater1317_in[12], zll_main_rotater1317_in[11], zll_main_rotater1317_in[10], zll_main_rotater1317_in[9], zll_main_rotater1317_in[8], zll_main_rotater1317_in[7], zll_main_rotater1317_in[6], zll_main_rotater1317_in[5], zll_main_rotater1317_in[4], zll_main_rotater1317_in[3], zll_main_rotater1317_in[2], zll_main_rotater1317_in[1], zll_main_rotater1317_in[0]};
  assign zll_main_rotater1319_in = {zll_main_rotater1321_in[31], zll_main_rotater1321_in[30], zll_main_rotater1321_in[25], zll_main_rotater1321_in[29], zll_main_rotater1321_in[28], zll_main_rotater1321_in[27], zll_main_rotater1321_in[26], zll_main_rotater1321_in[24], zll_main_rotater1321_in[23], zll_main_rotater1321_in[22], zll_main_rotater1321_in[21], zll_main_rotater1321_in[20], zll_main_rotater1321_in[19], zll_main_rotater1321_in[18], zll_main_rotater1321_in[17], zll_main_rotater1321_in[16], zll_main_rotater1321_in[15], zll_main_rotater1321_in[14], zll_main_rotater1321_in[13], zll_main_rotater1321_in[12], zll_main_rotater1321_in[11], zll_main_rotater1321_in[10], zll_main_rotater1321_in[9], zll_main_rotater1321_in[8], zll_main_rotater1321_in[7], zll_main_rotater1321_in[6], zll_main_rotater1321_in[5], zll_main_rotater1321_in[4], zll_main_rotater1321_in[3], zll_main_rotater1321_in[2], zll_main_rotater1321_in[1], zll_main_rotater1321_in[0]};
  assign zll_main_rotater1326_in = {zll_main_rotater1319_in[31], zll_main_rotater1319_in[30], zll_main_rotater1319_in[29], zll_main_rotater1319_in[24], zll_main_rotater1319_in[28], zll_main_rotater1319_in[27], zll_main_rotater1319_in[26], zll_main_rotater1319_in[25], zll_main_rotater1319_in[23], zll_main_rotater1319_in[22], zll_main_rotater1319_in[21], zll_main_rotater1319_in[20], zll_main_rotater1319_in[19], zll_main_rotater1319_in[18], zll_main_rotater1319_in[17], zll_main_rotater1319_in[16], zll_main_rotater1319_in[15], zll_main_rotater1319_in[14], zll_main_rotater1319_in[13], zll_main_rotater1319_in[12], zll_main_rotater1319_in[11], zll_main_rotater1319_in[10], zll_main_rotater1319_in[9], zll_main_rotater1319_in[8], zll_main_rotater1319_in[7], zll_main_rotater1319_in[6], zll_main_rotater1319_in[5], zll_main_rotater1319_in[4], zll_main_rotater1319_in[3], zll_main_rotater1319_in[2], zll_main_rotater1319_in[1], zll_main_rotater1319_in[0]};
  assign zll_main_rotater1331_in = {zll_main_rotater1326_in[31], zll_main_rotater1326_in[30], zll_main_rotater1326_in[29], zll_main_rotater1326_in[28], zll_main_rotater1326_in[27], zll_main_rotater1326_in[26], zll_main_rotater1326_in[25], zll_main_rotater1326_in[22], zll_main_rotater1326_in[24], zll_main_rotater1326_in[23], zll_main_rotater1326_in[21], zll_main_rotater1326_in[20], zll_main_rotater1326_in[19], zll_main_rotater1326_in[18], zll_main_rotater1326_in[17], zll_main_rotater1326_in[16], zll_main_rotater1326_in[15], zll_main_rotater1326_in[14], zll_main_rotater1326_in[13], zll_main_rotater1326_in[12], zll_main_rotater1326_in[11], zll_main_rotater1326_in[10], zll_main_rotater1326_in[9], zll_main_rotater1326_in[8], zll_main_rotater1326_in[7], zll_main_rotater1326_in[6], zll_main_rotater1326_in[5], zll_main_rotater1326_in[4], zll_main_rotater1326_in[3], zll_main_rotater1326_in[2], zll_main_rotater1326_in[1], zll_main_rotater1326_in[0]};
  assign zll_main_rotater1310_in = {zll_main_rotater1331_in[31], zll_main_rotater1331_in[30], zll_main_rotater1331_in[29], zll_main_rotater1331_in[28], zll_main_rotater1331_in[27], zll_main_rotater1331_in[26], zll_main_rotater1331_in[25], zll_main_rotater1331_in[24], zll_main_rotater1331_in[23], zll_main_rotater1331_in[21], zll_main_rotater1331_in[22], zll_main_rotater1331_in[20], zll_main_rotater1331_in[19], zll_main_rotater1331_in[18], zll_main_rotater1331_in[17], zll_main_rotater1331_in[16], zll_main_rotater1331_in[15], zll_main_rotater1331_in[14], zll_main_rotater1331_in[13], zll_main_rotater1331_in[12], zll_main_rotater1331_in[11], zll_main_rotater1331_in[10], zll_main_rotater1331_in[9], zll_main_rotater1331_in[8], zll_main_rotater1331_in[7], zll_main_rotater1331_in[6], zll_main_rotater1331_in[5], zll_main_rotater1331_in[4], zll_main_rotater1331_in[3], zll_main_rotater1331_in[2], zll_main_rotater1331_in[1], zll_main_rotater1331_in[0]};
  assign zll_main_rotater1311_in = {zll_main_rotater1310_in[20], zll_main_rotater1310_in[31], zll_main_rotater1310_in[30], zll_main_rotater1310_in[29], zll_main_rotater1310_in[28], zll_main_rotater1310_in[27], zll_main_rotater1310_in[26], zll_main_rotater1310_in[25], zll_main_rotater1310_in[24], zll_main_rotater1310_in[23], zll_main_rotater1310_in[22], zll_main_rotater1310_in[21], zll_main_rotater1310_in[19], zll_main_rotater1310_in[18], zll_main_rotater1310_in[17], zll_main_rotater1310_in[16], zll_main_rotater1310_in[15], zll_main_rotater1310_in[14], zll_main_rotater1310_in[13], zll_main_rotater1310_in[12], zll_main_rotater1310_in[11], zll_main_rotater1310_in[10], zll_main_rotater1310_in[9], zll_main_rotater1310_in[8], zll_main_rotater1310_in[7], zll_main_rotater1310_in[6], zll_main_rotater1310_in[5], zll_main_rotater1310_in[4], zll_main_rotater1310_in[3], zll_main_rotater1310_in[2], zll_main_rotater1310_in[1], zll_main_rotater1310_in[0]};
  assign zll_main_rotater131_in = {zll_main_rotater1311_in[31], zll_main_rotater1311_in[30], zll_main_rotater1311_in[29], zll_main_rotater1311_in[28], zll_main_rotater1311_in[27], zll_main_rotater1311_in[26], zll_main_rotater1311_in[25], zll_main_rotater1311_in[24], zll_main_rotater1311_in[23], zll_main_rotater1311_in[22], zll_main_rotater1311_in[19], zll_main_rotater1311_in[21], zll_main_rotater1311_in[20], zll_main_rotater1311_in[18], zll_main_rotater1311_in[17], zll_main_rotater1311_in[16], zll_main_rotater1311_in[15], zll_main_rotater1311_in[14], zll_main_rotater1311_in[13], zll_main_rotater1311_in[12], zll_main_rotater1311_in[11], zll_main_rotater1311_in[10], zll_main_rotater1311_in[9], zll_main_rotater1311_in[8], zll_main_rotater1311_in[7], zll_main_rotater1311_in[6], zll_main_rotater1311_in[5], zll_main_rotater1311_in[4], zll_main_rotater1311_in[3], zll_main_rotater1311_in[2], zll_main_rotater1311_in[1], zll_main_rotater1311_in[0]};
  assign zll_main_rotater1325_in = {zll_main_rotater131_in[31], zll_main_rotater131_in[30], zll_main_rotater131_in[29], zll_main_rotater131_in[28], zll_main_rotater131_in[27], zll_main_rotater131_in[26], zll_main_rotater131_in[25], zll_main_rotater131_in[24], zll_main_rotater131_in[23], zll_main_rotater131_in[18], zll_main_rotater131_in[22], zll_main_rotater131_in[21], zll_main_rotater131_in[20], zll_main_rotater131_in[19], zll_main_rotater131_in[17], zll_main_rotater131_in[16], zll_main_rotater131_in[15], zll_main_rotater131_in[14], zll_main_rotater131_in[13], zll_main_rotater131_in[12], zll_main_rotater131_in[11], zll_main_rotater131_in[10], zll_main_rotater131_in[9], zll_main_rotater131_in[8], zll_main_rotater131_in[7], zll_main_rotater131_in[6], zll_main_rotater131_in[5], zll_main_rotater131_in[4], zll_main_rotater131_in[3], zll_main_rotater131_in[2], zll_main_rotater131_in[1], zll_main_rotater131_in[0]};
  assign zll_main_rotater1329_in = {zll_main_rotater1325_in[31], zll_main_rotater1325_in[30], zll_main_rotater1325_in[29], zll_main_rotater1325_in[28], zll_main_rotater1325_in[27], zll_main_rotater1325_in[26], zll_main_rotater1325_in[25], zll_main_rotater1325_in[24], zll_main_rotater1325_in[23], zll_main_rotater1325_in[22], zll_main_rotater1325_in[21], zll_main_rotater1325_in[20], zll_main_rotater1325_in[19], zll_main_rotater1325_in[17], zll_main_rotater1325_in[18], zll_main_rotater1325_in[16], zll_main_rotater1325_in[15], zll_main_rotater1325_in[14], zll_main_rotater1325_in[13], zll_main_rotater1325_in[12], zll_main_rotater1325_in[11], zll_main_rotater1325_in[10], zll_main_rotater1325_in[9], zll_main_rotater1325_in[8], zll_main_rotater1325_in[7], zll_main_rotater1325_in[6], zll_main_rotater1325_in[5], zll_main_rotater1325_in[4], zll_main_rotater1325_in[3], zll_main_rotater1325_in[2], zll_main_rotater1325_in[1], zll_main_rotater1325_in[0]};
  assign zll_main_rotater1312_in = {zll_main_rotater1329_in[31], zll_main_rotater1329_in[30], zll_main_rotater1329_in[29], zll_main_rotater1329_in[28], zll_main_rotater1329_in[27], zll_main_rotater1329_in[26], zll_main_rotater1329_in[25], zll_main_rotater1329_in[16], zll_main_rotater1329_in[24], zll_main_rotater1329_in[23], zll_main_rotater1329_in[22], zll_main_rotater1329_in[21], zll_main_rotater1329_in[20], zll_main_rotater1329_in[19], zll_main_rotater1329_in[18], zll_main_rotater1329_in[17], zll_main_rotater1329_in[15], zll_main_rotater1329_in[14], zll_main_rotater1329_in[13], zll_main_rotater1329_in[12], zll_main_rotater1329_in[11], zll_main_rotater1329_in[10], zll_main_rotater1329_in[9], zll_main_rotater1329_in[8], zll_main_rotater1329_in[7], zll_main_rotater1329_in[6], zll_main_rotater1329_in[5], zll_main_rotater1329_in[4], zll_main_rotater1329_in[3], zll_main_rotater1329_in[2], zll_main_rotater1329_in[1], zll_main_rotater1329_in[0]};
  assign zll_main_rotater132_in = {zll_main_rotater1312_in[31], zll_main_rotater1312_in[30], zll_main_rotater1312_in[29], zll_main_rotater1312_in[28], zll_main_rotater1312_in[27], zll_main_rotater1312_in[26], zll_main_rotater1312_in[25], zll_main_rotater1312_in[15], zll_main_rotater1312_in[24], zll_main_rotater1312_in[23], zll_main_rotater1312_in[22], zll_main_rotater1312_in[21], zll_main_rotater1312_in[20], zll_main_rotater1312_in[19], zll_main_rotater1312_in[18], zll_main_rotater1312_in[17], zll_main_rotater1312_in[16], zll_main_rotater1312_in[14], zll_main_rotater1312_in[13], zll_main_rotater1312_in[12], zll_main_rotater1312_in[11], zll_main_rotater1312_in[10], zll_main_rotater1312_in[9], zll_main_rotater1312_in[8], zll_main_rotater1312_in[7], zll_main_rotater1312_in[6], zll_main_rotater1312_in[5], zll_main_rotater1312_in[4], zll_main_rotater1312_in[3], zll_main_rotater1312_in[2], zll_main_rotater1312_in[1], zll_main_rotater1312_in[0]};
  assign zll_main_rotater1327_in = {zll_main_rotater132_in[31], zll_main_rotater132_in[30], zll_main_rotater132_in[29], zll_main_rotater132_in[28], zll_main_rotater132_in[27], zll_main_rotater132_in[26], zll_main_rotater132_in[25], zll_main_rotater132_in[24], zll_main_rotater132_in[23], zll_main_rotater132_in[22], zll_main_rotater132_in[21], zll_main_rotater132_in[20], zll_main_rotater132_in[14], zll_main_rotater132_in[19], zll_main_rotater132_in[18], zll_main_rotater132_in[17], zll_main_rotater132_in[16], zll_main_rotater132_in[15], zll_main_rotater132_in[13], zll_main_rotater132_in[12], zll_main_rotater132_in[11], zll_main_rotater132_in[10], zll_main_rotater132_in[9], zll_main_rotater132_in[8], zll_main_rotater132_in[7], zll_main_rotater132_in[6], zll_main_rotater132_in[5], zll_main_rotater132_in[4], zll_main_rotater132_in[3], zll_main_rotater132_in[2], zll_main_rotater132_in[1], zll_main_rotater132_in[0]};
  assign zll_main_rotater1322_in = {zll_main_rotater1327_in[31], zll_main_rotater1327_in[30], zll_main_rotater1327_in[29], zll_main_rotater1327_in[28], zll_main_rotater1327_in[27], zll_main_rotater1327_in[26], zll_main_rotater1327_in[25], zll_main_rotater1327_in[24], zll_main_rotater1327_in[23], zll_main_rotater1327_in[22], zll_main_rotater1327_in[21], zll_main_rotater1327_in[20], zll_main_rotater1327_in[13], zll_main_rotater1327_in[19], zll_main_rotater1327_in[18], zll_main_rotater1327_in[17], zll_main_rotater1327_in[16], zll_main_rotater1327_in[15], zll_main_rotater1327_in[14], zll_main_rotater1327_in[12], zll_main_rotater1327_in[11], zll_main_rotater1327_in[10], zll_main_rotater1327_in[9], zll_main_rotater1327_in[8], zll_main_rotater1327_in[7], zll_main_rotater1327_in[6], zll_main_rotater1327_in[5], zll_main_rotater1327_in[4], zll_main_rotater1327_in[3], zll_main_rotater1327_in[2], zll_main_rotater1327_in[1], zll_main_rotater1327_in[0]};
  assign zll_main_rotater137_in = {zll_main_rotater1322_in[31], zll_main_rotater1322_in[30], zll_main_rotater1322_in[29], zll_main_rotater1322_in[28], zll_main_rotater1322_in[27], zll_main_rotater1322_in[26], zll_main_rotater1322_in[25], zll_main_rotater1322_in[24], zll_main_rotater1322_in[23], zll_main_rotater1322_in[22], zll_main_rotater1322_in[21], zll_main_rotater1322_in[20], zll_main_rotater1322_in[19], zll_main_rotater1322_in[18], zll_main_rotater1322_in[17], zll_main_rotater1322_in[16], zll_main_rotater1322_in[12], zll_main_rotater1322_in[15], zll_main_rotater1322_in[14], zll_main_rotater1322_in[13], zll_main_rotater1322_in[11], zll_main_rotater1322_in[10], zll_main_rotater1322_in[9], zll_main_rotater1322_in[8], zll_main_rotater1322_in[7], zll_main_rotater1322_in[6], zll_main_rotater1322_in[5], zll_main_rotater1322_in[4], zll_main_rotater1322_in[3], zll_main_rotater1322_in[2], zll_main_rotater1322_in[1], zll_main_rotater1322_in[0]};
  assign zll_main_rotater134_in = {zll_main_rotater137_in[31], zll_main_rotater137_in[30], zll_main_rotater137_in[29], zll_main_rotater137_in[28], zll_main_rotater137_in[11], zll_main_rotater137_in[27], zll_main_rotater137_in[26], zll_main_rotater137_in[25], zll_main_rotater137_in[24], zll_main_rotater137_in[23], zll_main_rotater137_in[22], zll_main_rotater137_in[21], zll_main_rotater137_in[20], zll_main_rotater137_in[19], zll_main_rotater137_in[18], zll_main_rotater137_in[17], zll_main_rotater137_in[16], zll_main_rotater137_in[15], zll_main_rotater137_in[14], zll_main_rotater137_in[13], zll_main_rotater137_in[12], zll_main_rotater137_in[10], zll_main_rotater137_in[9], zll_main_rotater137_in[8], zll_main_rotater137_in[7], zll_main_rotater137_in[6], zll_main_rotater137_in[5], zll_main_rotater137_in[4], zll_main_rotater137_in[3], zll_main_rotater137_in[2], zll_main_rotater137_in[1], zll_main_rotater137_in[0]};
  assign zll_main_rotater1330_in = {zll_main_rotater134_in[31], zll_main_rotater134_in[30], zll_main_rotater134_in[29], zll_main_rotater134_in[28], zll_main_rotater134_in[27], zll_main_rotater134_in[26], zll_main_rotater134_in[25], zll_main_rotater134_in[24], zll_main_rotater134_in[23], zll_main_rotater134_in[22], zll_main_rotater134_in[21], zll_main_rotater134_in[20], zll_main_rotater134_in[19], zll_main_rotater134_in[18], zll_main_rotater134_in[17], zll_main_rotater134_in[16], zll_main_rotater134_in[15], zll_main_rotater134_in[14], zll_main_rotater134_in[10], zll_main_rotater134_in[13], zll_main_rotater134_in[12], zll_main_rotater134_in[11], zll_main_rotater134_in[9], zll_main_rotater134_in[8], zll_main_rotater134_in[7], zll_main_rotater134_in[6], zll_main_rotater134_in[5], zll_main_rotater134_in[4], zll_main_rotater134_in[3], zll_main_rotater134_in[2], zll_main_rotater134_in[1], zll_main_rotater134_in[0]};
  assign zll_main_rotater1320_in = {zll_main_rotater1330_in[31], zll_main_rotater1330_in[30], zll_main_rotater1330_in[29], zll_main_rotater1330_in[28], zll_main_rotater1330_in[27], zll_main_rotater1330_in[26], zll_main_rotater1330_in[25], zll_main_rotater1330_in[24], zll_main_rotater1330_in[23], zll_main_rotater1330_in[9], zll_main_rotater1330_in[22], zll_main_rotater1330_in[21], zll_main_rotater1330_in[20], zll_main_rotater1330_in[19], zll_main_rotater1330_in[18], zll_main_rotater1330_in[17], zll_main_rotater1330_in[16], zll_main_rotater1330_in[15], zll_main_rotater1330_in[14], zll_main_rotater1330_in[13], zll_main_rotater1330_in[12], zll_main_rotater1330_in[11], zll_main_rotater1330_in[10], zll_main_rotater1330_in[8], zll_main_rotater1330_in[7], zll_main_rotater1330_in[6], zll_main_rotater1330_in[5], zll_main_rotater1330_in[4], zll_main_rotater1330_in[3], zll_main_rotater1330_in[2], zll_main_rotater1330_in[1], zll_main_rotater1330_in[0]};
  assign zll_main_rotater1315_in = {zll_main_rotater1320_in[31], zll_main_rotater1320_in[30], zll_main_rotater1320_in[29], zll_main_rotater1320_in[28], zll_main_rotater1320_in[27], zll_main_rotater1320_in[26], zll_main_rotater1320_in[25], zll_main_rotater1320_in[24], zll_main_rotater1320_in[23], zll_main_rotater1320_in[22], zll_main_rotater1320_in[21], zll_main_rotater1320_in[20], zll_main_rotater1320_in[19], zll_main_rotater1320_in[18], zll_main_rotater1320_in[17], zll_main_rotater1320_in[16], zll_main_rotater1320_in[15], zll_main_rotater1320_in[14], zll_main_rotater1320_in[13], zll_main_rotater1320_in[12], zll_main_rotater1320_in[11], zll_main_rotater1320_in[10], zll_main_rotater1320_in[8], zll_main_rotater1320_in[9], zll_main_rotater1320_in[7], zll_main_rotater1320_in[6], zll_main_rotater1320_in[5], zll_main_rotater1320_in[4], zll_main_rotater1320_in[3], zll_main_rotater1320_in[2], zll_main_rotater1320_in[1], zll_main_rotater1320_in[0]};
  assign zll_main_rotater1313_in = {zll_main_rotater1315_in[31], zll_main_rotater1315_in[30], zll_main_rotater1315_in[29], zll_main_rotater1315_in[28], zll_main_rotater1315_in[27], zll_main_rotater1315_in[7], zll_main_rotater1315_in[26], zll_main_rotater1315_in[25], zll_main_rotater1315_in[24], zll_main_rotater1315_in[23], zll_main_rotater1315_in[22], zll_main_rotater1315_in[21], zll_main_rotater1315_in[20], zll_main_rotater1315_in[19], zll_main_rotater1315_in[18], zll_main_rotater1315_in[17], zll_main_rotater1315_in[16], zll_main_rotater1315_in[15], zll_main_rotater1315_in[14], zll_main_rotater1315_in[13], zll_main_rotater1315_in[12], zll_main_rotater1315_in[11], zll_main_rotater1315_in[10], zll_main_rotater1315_in[9], zll_main_rotater1315_in[8], zll_main_rotater1315_in[6], zll_main_rotater1315_in[5], zll_main_rotater1315_in[4], zll_main_rotater1315_in[3], zll_main_rotater1315_in[2], zll_main_rotater1315_in[1], zll_main_rotater1315_in[0]};
  assign zll_main_rotater13_in = {zll_main_rotater1313_in[31], zll_main_rotater1313_in[30], zll_main_rotater1313_in[29], zll_main_rotater1313_in[28], zll_main_rotater1313_in[27], zll_main_rotater1313_in[26], zll_main_rotater1313_in[25], zll_main_rotater1313_in[6], zll_main_rotater1313_in[24], zll_main_rotater1313_in[23], zll_main_rotater1313_in[22], zll_main_rotater1313_in[21], zll_main_rotater1313_in[20], zll_main_rotater1313_in[19], zll_main_rotater1313_in[18], zll_main_rotater1313_in[17], zll_main_rotater1313_in[16], zll_main_rotater1313_in[15], zll_main_rotater1313_in[14], zll_main_rotater1313_in[13], zll_main_rotater1313_in[12], zll_main_rotater1313_in[11], zll_main_rotater1313_in[10], zll_main_rotater1313_in[9], zll_main_rotater1313_in[8], zll_main_rotater1313_in[7], zll_main_rotater1313_in[5], zll_main_rotater1313_in[4], zll_main_rotater1313_in[3], zll_main_rotater1313_in[2], zll_main_rotater1313_in[1], zll_main_rotater1313_in[0]};
  assign zll_main_rotater136_in = {zll_main_rotater13_in[31], zll_main_rotater13_in[5], zll_main_rotater13_in[30], zll_main_rotater13_in[29], zll_main_rotater13_in[28], zll_main_rotater13_in[27], zll_main_rotater13_in[26], zll_main_rotater13_in[25], zll_main_rotater13_in[24], zll_main_rotater13_in[23], zll_main_rotater13_in[22], zll_main_rotater13_in[21], zll_main_rotater13_in[20], zll_main_rotater13_in[19], zll_main_rotater13_in[18], zll_main_rotater13_in[17], zll_main_rotater13_in[16], zll_main_rotater13_in[15], zll_main_rotater13_in[14], zll_main_rotater13_in[13], zll_main_rotater13_in[12], zll_main_rotater13_in[11], zll_main_rotater13_in[10], zll_main_rotater13_in[9], zll_main_rotater13_in[8], zll_main_rotater13_in[7], zll_main_rotater13_in[6], zll_main_rotater13_in[4], zll_main_rotater13_in[3], zll_main_rotater13_in[2], zll_main_rotater13_in[1], zll_main_rotater13_in[0]};
  assign zll_main_rotater1318_in = {zll_main_rotater136_in[31], zll_main_rotater136_in[30], zll_main_rotater136_in[29], zll_main_rotater136_in[28], zll_main_rotater136_in[27], zll_main_rotater136_in[26], zll_main_rotater136_in[25], zll_main_rotater136_in[24], zll_main_rotater136_in[23], zll_main_rotater136_in[22], zll_main_rotater136_in[21], zll_main_rotater136_in[20], zll_main_rotater136_in[19], zll_main_rotater136_in[18], zll_main_rotater136_in[17], zll_main_rotater136_in[16], zll_main_rotater136_in[15], zll_main_rotater136_in[4], zll_main_rotater136_in[14], zll_main_rotater136_in[13], zll_main_rotater136_in[12], zll_main_rotater136_in[11], zll_main_rotater136_in[10], zll_main_rotater136_in[9], zll_main_rotater136_in[8], zll_main_rotater136_in[7], zll_main_rotater136_in[6], zll_main_rotater136_in[5], zll_main_rotater136_in[3], zll_main_rotater136_in[2], zll_main_rotater136_in[1], zll_main_rotater136_in[0]};
  assign zll_main_rotater135_in = {zll_main_rotater1318_in[31], zll_main_rotater1318_in[30], zll_main_rotater1318_in[29], zll_main_rotater1318_in[28], zll_main_rotater1318_in[27], zll_main_rotater1318_in[26], zll_main_rotater1318_in[25], zll_main_rotater1318_in[24], zll_main_rotater1318_in[23], zll_main_rotater1318_in[22], zll_main_rotater1318_in[21], zll_main_rotater1318_in[20], zll_main_rotater1318_in[19], zll_main_rotater1318_in[18], zll_main_rotater1318_in[17], zll_main_rotater1318_in[3], zll_main_rotater1318_in[16], zll_main_rotater1318_in[15], zll_main_rotater1318_in[14], zll_main_rotater1318_in[13], zll_main_rotater1318_in[12], zll_main_rotater1318_in[11], zll_main_rotater1318_in[10], zll_main_rotater1318_in[9], zll_main_rotater1318_in[8], zll_main_rotater1318_in[7], zll_main_rotater1318_in[6], zll_main_rotater1318_in[5], zll_main_rotater1318_in[4], zll_main_rotater1318_in[2], zll_main_rotater1318_in[1], zll_main_rotater1318_in[0]};
  assign zll_main_rotater133_in = {zll_main_rotater135_in[31], zll_main_rotater135_in[2], zll_main_rotater135_in[30], zll_main_rotater135_in[29], zll_main_rotater135_in[28], zll_main_rotater135_in[27], zll_main_rotater135_in[26], zll_main_rotater135_in[25], zll_main_rotater135_in[24], zll_main_rotater135_in[23], zll_main_rotater135_in[22], zll_main_rotater135_in[21], zll_main_rotater135_in[20], zll_main_rotater135_in[19], zll_main_rotater135_in[18], zll_main_rotater135_in[17], zll_main_rotater135_in[16], zll_main_rotater135_in[15], zll_main_rotater135_in[14], zll_main_rotater135_in[13], zll_main_rotater135_in[12], zll_main_rotater135_in[11], zll_main_rotater135_in[10], zll_main_rotater135_in[9], zll_main_rotater135_in[8], zll_main_rotater135_in[7], zll_main_rotater135_in[6], zll_main_rotater135_in[5], zll_main_rotater135_in[4], zll_main_rotater135_in[3], zll_main_rotater135_in[1], zll_main_rotater135_in[0]};
  assign zll_main_rotater1314_in = {zll_main_rotater133_in[31], zll_main_rotater133_in[30], zll_main_rotater133_in[29], zll_main_rotater133_in[28], zll_main_rotater133_in[27], zll_main_rotater133_in[26], zll_main_rotater133_in[1], zll_main_rotater133_in[25], zll_main_rotater133_in[24], zll_main_rotater133_in[23], zll_main_rotater133_in[22], zll_main_rotater133_in[21], zll_main_rotater133_in[20], zll_main_rotater133_in[19], zll_main_rotater133_in[18], zll_main_rotater133_in[17], zll_main_rotater133_in[16], zll_main_rotater133_in[15], zll_main_rotater133_in[14], zll_main_rotater133_in[13], zll_main_rotater133_in[12], zll_main_rotater133_in[11], zll_main_rotater133_in[10], zll_main_rotater133_in[9], zll_main_rotater133_in[8], zll_main_rotater133_in[7], zll_main_rotater133_in[6], zll_main_rotater133_in[5], zll_main_rotater133_in[4], zll_main_rotater133_in[3], zll_main_rotater133_in[2], zll_main_rotater133_in[0]};
  assign xorw32_inR4 = {{zll_main_rotater237_in[27], zll_main_rotater237_in[0], zll_main_rotater237_in[8], zll_main_rotater237_in[18], zll_main_rotater237_in[11], zll_main_rotater237_in[3], zll_main_rotater237_in[17], zll_main_rotater237_in[28], zll_main_rotater237_in[22], zll_main_rotater237_in[10], zll_main_rotater237_in[14], zll_main_rotater237_in[13], zll_main_rotater237_in[31], zll_main_rotater237_in[25], zll_main_rotater237_in[16], zll_main_rotater237_in[29], zll_main_rotater237_in[24], zll_main_rotater237_in[9], zll_main_rotater237_in[26], zll_main_rotater237_in[21], zll_main_rotater237_in[1], zll_main_rotater237_in[19], zll_main_rotater237_in[4], zll_main_rotater237_in[12], zll_main_rotater237_in[5], zll_main_rotater237_in[6], zll_main_rotater237_in[20], zll_main_rotater237_in[30], zll_main_rotater237_in[23], zll_main_rotater237_in[2], zll_main_rotater237_in[7], zll_main_rotater237_in[15]}, {zll_main_rotater1314_in[6], zll_main_rotater1314_in[24], zll_main_rotater1314_in[5], zll_main_rotater1314_in[17], zll_main_rotater1314_in[2], zll_main_rotater1314_in[23], zll_main_rotater1314_in[21], zll_main_rotater1314_in[29], zll_main_rotater1314_in[11], zll_main_rotater1314_in[14], zll_main_rotater1314_in[30], zll_main_rotater1314_in[25], zll_main_rotater1314_in[0], zll_main_rotater1314_in[27], zll_main_rotater1314_in[8], zll_main_rotater1314_in[28], zll_main_rotater1314_in[20], zll_main_rotater1314_in[19], zll_main_rotater1314_in[15], zll_main_rotater1314_in[26], zll_main_rotater1314_in[22], zll_main_rotater1314_in[1], zll_main_rotater1314_in[13], zll_main_rotater1314_in[4], zll_main_rotater1314_in[31], zll_main_rotater1314_in[7], zll_main_rotater1314_in[12], zll_main_rotater1314_in[3], zll_main_rotater1314_in[16], zll_main_rotater1314_in[18], zll_main_rotater1314_in[9], zll_main_rotater1314_in[10]}};
  xorW32  instR13 (xorw32_inR4[63:32], xorw32_inR4[31:0], extresR11[31:0]);
  assign main_rotater22_in = main_bigsigma0_in[31:0];
  assign zll_main_rotater227_in = main_rotater22_in[31:0];
  assign zll_main_rotater2213_in = {zll_main_rotater227_in[29], zll_main_rotater227_in[31], zll_main_rotater227_in[30], zll_main_rotater227_in[28], zll_main_rotater227_in[27], zll_main_rotater227_in[26], zll_main_rotater227_in[25], zll_main_rotater227_in[24], zll_main_rotater227_in[23], zll_main_rotater227_in[22], zll_main_rotater227_in[21], zll_main_rotater227_in[20], zll_main_rotater227_in[19], zll_main_rotater227_in[18], zll_main_rotater227_in[17], zll_main_rotater227_in[16], zll_main_rotater227_in[15], zll_main_rotater227_in[14], zll_main_rotater227_in[13], zll_main_rotater227_in[12], zll_main_rotater227_in[11], zll_main_rotater227_in[10], zll_main_rotater227_in[9], zll_main_rotater227_in[8], zll_main_rotater227_in[7], zll_main_rotater227_in[6], zll_main_rotater227_in[5], zll_main_rotater227_in[4], zll_main_rotater227_in[3], zll_main_rotater227_in[2], zll_main_rotater227_in[1], zll_main_rotater227_in[0]};
  assign zll_main_rotater2229_in = {zll_main_rotater2213_in[28], zll_main_rotater2213_in[31], zll_main_rotater2213_in[30], zll_main_rotater2213_in[29], zll_main_rotater2213_in[27], zll_main_rotater2213_in[26], zll_main_rotater2213_in[25], zll_main_rotater2213_in[24], zll_main_rotater2213_in[23], zll_main_rotater2213_in[22], zll_main_rotater2213_in[21], zll_main_rotater2213_in[20], zll_main_rotater2213_in[19], zll_main_rotater2213_in[18], zll_main_rotater2213_in[17], zll_main_rotater2213_in[16], zll_main_rotater2213_in[15], zll_main_rotater2213_in[14], zll_main_rotater2213_in[13], zll_main_rotater2213_in[12], zll_main_rotater2213_in[11], zll_main_rotater2213_in[10], zll_main_rotater2213_in[9], zll_main_rotater2213_in[8], zll_main_rotater2213_in[7], zll_main_rotater2213_in[6], zll_main_rotater2213_in[5], zll_main_rotater2213_in[4], zll_main_rotater2213_in[3], zll_main_rotater2213_in[2], zll_main_rotater2213_in[1], zll_main_rotater2213_in[0]};
  assign zll_main_rotater2230_in = {zll_main_rotater2229_in[31], zll_main_rotater2229_in[30], zll_main_rotater2229_in[27], zll_main_rotater2229_in[29], zll_main_rotater2229_in[28], zll_main_rotater2229_in[26], zll_main_rotater2229_in[25], zll_main_rotater2229_in[24], zll_main_rotater2229_in[23], zll_main_rotater2229_in[22], zll_main_rotater2229_in[21], zll_main_rotater2229_in[20], zll_main_rotater2229_in[19], zll_main_rotater2229_in[18], zll_main_rotater2229_in[17], zll_main_rotater2229_in[16], zll_main_rotater2229_in[15], zll_main_rotater2229_in[14], zll_main_rotater2229_in[13], zll_main_rotater2229_in[12], zll_main_rotater2229_in[11], zll_main_rotater2229_in[10], zll_main_rotater2229_in[9], zll_main_rotater2229_in[8], zll_main_rotater2229_in[7], zll_main_rotater2229_in[6], zll_main_rotater2229_in[5], zll_main_rotater2229_in[4], zll_main_rotater2229_in[3], zll_main_rotater2229_in[2], zll_main_rotater2229_in[1], zll_main_rotater2229_in[0]};
  assign zll_main_rotater2214_in = {zll_main_rotater2230_in[31], zll_main_rotater2230_in[30], zll_main_rotater2230_in[29], zll_main_rotater2230_in[25], zll_main_rotater2230_in[28], zll_main_rotater2230_in[27], zll_main_rotater2230_in[26], zll_main_rotater2230_in[24], zll_main_rotater2230_in[23], zll_main_rotater2230_in[22], zll_main_rotater2230_in[21], zll_main_rotater2230_in[20], zll_main_rotater2230_in[19], zll_main_rotater2230_in[18], zll_main_rotater2230_in[17], zll_main_rotater2230_in[16], zll_main_rotater2230_in[15], zll_main_rotater2230_in[14], zll_main_rotater2230_in[13], zll_main_rotater2230_in[12], zll_main_rotater2230_in[11], zll_main_rotater2230_in[10], zll_main_rotater2230_in[9], zll_main_rotater2230_in[8], zll_main_rotater2230_in[7], zll_main_rotater2230_in[6], zll_main_rotater2230_in[5], zll_main_rotater2230_in[4], zll_main_rotater2230_in[3], zll_main_rotater2230_in[2], zll_main_rotater2230_in[1], zll_main_rotater2230_in[0]};
  assign zll_main_rotater2226_in = {zll_main_rotater2214_in[31], zll_main_rotater2214_in[24], zll_main_rotater2214_in[30], zll_main_rotater2214_in[29], zll_main_rotater2214_in[28], zll_main_rotater2214_in[27], zll_main_rotater2214_in[26], zll_main_rotater2214_in[25], zll_main_rotater2214_in[23], zll_main_rotater2214_in[22], zll_main_rotater2214_in[21], zll_main_rotater2214_in[20], zll_main_rotater2214_in[19], zll_main_rotater2214_in[18], zll_main_rotater2214_in[17], zll_main_rotater2214_in[16], zll_main_rotater2214_in[15], zll_main_rotater2214_in[14], zll_main_rotater2214_in[13], zll_main_rotater2214_in[12], zll_main_rotater2214_in[11], zll_main_rotater2214_in[10], zll_main_rotater2214_in[9], zll_main_rotater2214_in[8], zll_main_rotater2214_in[7], zll_main_rotater2214_in[6], zll_main_rotater2214_in[5], zll_main_rotater2214_in[4], zll_main_rotater2214_in[3], zll_main_rotater2214_in[2], zll_main_rotater2214_in[1], zll_main_rotater2214_in[0]};
  assign zll_main_rotater2228_in = {zll_main_rotater2226_in[31], zll_main_rotater2226_in[30], zll_main_rotater2226_in[29], zll_main_rotater2226_in[28], zll_main_rotater2226_in[27], zll_main_rotater2226_in[26], zll_main_rotater2226_in[25], zll_main_rotater2226_in[23], zll_main_rotater2226_in[24], zll_main_rotater2226_in[22], zll_main_rotater2226_in[21], zll_main_rotater2226_in[20], zll_main_rotater2226_in[19], zll_main_rotater2226_in[18], zll_main_rotater2226_in[17], zll_main_rotater2226_in[16], zll_main_rotater2226_in[15], zll_main_rotater2226_in[14], zll_main_rotater2226_in[13], zll_main_rotater2226_in[12], zll_main_rotater2226_in[11], zll_main_rotater2226_in[10], zll_main_rotater2226_in[9], zll_main_rotater2226_in[8], zll_main_rotater2226_in[7], zll_main_rotater2226_in[6], zll_main_rotater2226_in[5], zll_main_rotater2226_in[4], zll_main_rotater2226_in[3], zll_main_rotater2226_in[2], zll_main_rotater2226_in[1], zll_main_rotater2226_in[0]};
  assign zll_main_rotater221_in = {zll_main_rotater2228_in[31], zll_main_rotater2228_in[30], zll_main_rotater2228_in[29], zll_main_rotater2228_in[28], zll_main_rotater2228_in[27], zll_main_rotater2228_in[22], zll_main_rotater2228_in[26], zll_main_rotater2228_in[25], zll_main_rotater2228_in[24], zll_main_rotater2228_in[23], zll_main_rotater2228_in[21], zll_main_rotater2228_in[20], zll_main_rotater2228_in[19], zll_main_rotater2228_in[18], zll_main_rotater2228_in[17], zll_main_rotater2228_in[16], zll_main_rotater2228_in[15], zll_main_rotater2228_in[14], zll_main_rotater2228_in[13], zll_main_rotater2228_in[12], zll_main_rotater2228_in[11], zll_main_rotater2228_in[10], zll_main_rotater2228_in[9], zll_main_rotater2228_in[8], zll_main_rotater2228_in[7], zll_main_rotater2228_in[6], zll_main_rotater2228_in[5], zll_main_rotater2228_in[4], zll_main_rotater2228_in[3], zll_main_rotater2228_in[2], zll_main_rotater2228_in[1], zll_main_rotater2228_in[0]};
  assign zll_main_rotater2224_in = {zll_main_rotater221_in[31], zll_main_rotater221_in[30], zll_main_rotater221_in[29], zll_main_rotater221_in[21], zll_main_rotater221_in[28], zll_main_rotater221_in[27], zll_main_rotater221_in[26], zll_main_rotater221_in[25], zll_main_rotater221_in[24], zll_main_rotater221_in[23], zll_main_rotater221_in[22], zll_main_rotater221_in[20], zll_main_rotater221_in[19], zll_main_rotater221_in[18], zll_main_rotater221_in[17], zll_main_rotater221_in[16], zll_main_rotater221_in[15], zll_main_rotater221_in[14], zll_main_rotater221_in[13], zll_main_rotater221_in[12], zll_main_rotater221_in[11], zll_main_rotater221_in[10], zll_main_rotater221_in[9], zll_main_rotater221_in[8], zll_main_rotater221_in[7], zll_main_rotater221_in[6], zll_main_rotater221_in[5], zll_main_rotater221_in[4], zll_main_rotater221_in[3], zll_main_rotater221_in[2], zll_main_rotater221_in[1], zll_main_rotater221_in[0]};
  assign zll_main_rotater2211_in = {zll_main_rotater2224_in[31], zll_main_rotater2224_in[30], zll_main_rotater2224_in[29], zll_main_rotater2224_in[28], zll_main_rotater2224_in[27], zll_main_rotater2224_in[26], zll_main_rotater2224_in[25], zll_main_rotater2224_in[24], zll_main_rotater2224_in[23], zll_main_rotater2224_in[20], zll_main_rotater2224_in[22], zll_main_rotater2224_in[21], zll_main_rotater2224_in[19], zll_main_rotater2224_in[18], zll_main_rotater2224_in[17], zll_main_rotater2224_in[16], zll_main_rotater2224_in[15], zll_main_rotater2224_in[14], zll_main_rotater2224_in[13], zll_main_rotater2224_in[12], zll_main_rotater2224_in[11], zll_main_rotater2224_in[10], zll_main_rotater2224_in[9], zll_main_rotater2224_in[8], zll_main_rotater2224_in[7], zll_main_rotater2224_in[6], zll_main_rotater2224_in[5], zll_main_rotater2224_in[4], zll_main_rotater2224_in[3], zll_main_rotater2224_in[2], zll_main_rotater2224_in[1], zll_main_rotater2224_in[0]};
  assign zll_main_rotater224_in = {zll_main_rotater2211_in[31], zll_main_rotater2211_in[30], zll_main_rotater2211_in[29], zll_main_rotater2211_in[19], zll_main_rotater2211_in[28], zll_main_rotater2211_in[27], zll_main_rotater2211_in[26], zll_main_rotater2211_in[25], zll_main_rotater2211_in[24], zll_main_rotater2211_in[23], zll_main_rotater2211_in[22], zll_main_rotater2211_in[21], zll_main_rotater2211_in[20], zll_main_rotater2211_in[18], zll_main_rotater2211_in[17], zll_main_rotater2211_in[16], zll_main_rotater2211_in[15], zll_main_rotater2211_in[14], zll_main_rotater2211_in[13], zll_main_rotater2211_in[12], zll_main_rotater2211_in[11], zll_main_rotater2211_in[10], zll_main_rotater2211_in[9], zll_main_rotater2211_in[8], zll_main_rotater2211_in[7], zll_main_rotater2211_in[6], zll_main_rotater2211_in[5], zll_main_rotater2211_in[4], zll_main_rotater2211_in[3], zll_main_rotater2211_in[2], zll_main_rotater2211_in[1], zll_main_rotater2211_in[0]};
  assign zll_main_rotater2219_in = {zll_main_rotater224_in[31], zll_main_rotater224_in[30], zll_main_rotater224_in[29], zll_main_rotater224_in[28], zll_main_rotater224_in[27], zll_main_rotater224_in[18], zll_main_rotater224_in[26], zll_main_rotater224_in[25], zll_main_rotater224_in[24], zll_main_rotater224_in[23], zll_main_rotater224_in[22], zll_main_rotater224_in[21], zll_main_rotater224_in[20], zll_main_rotater224_in[19], zll_main_rotater224_in[17], zll_main_rotater224_in[16], zll_main_rotater224_in[15], zll_main_rotater224_in[14], zll_main_rotater224_in[13], zll_main_rotater224_in[12], zll_main_rotater224_in[11], zll_main_rotater224_in[10], zll_main_rotater224_in[9], zll_main_rotater224_in[8], zll_main_rotater224_in[7], zll_main_rotater224_in[6], zll_main_rotater224_in[5], zll_main_rotater224_in[4], zll_main_rotater224_in[3], zll_main_rotater224_in[2], zll_main_rotater224_in[1], zll_main_rotater224_in[0]};
  assign zll_main_rotater2222_in = {zll_main_rotater2219_in[31], zll_main_rotater2219_in[30], zll_main_rotater2219_in[29], zll_main_rotater2219_in[28], zll_main_rotater2219_in[27], zll_main_rotater2219_in[26], zll_main_rotater2219_in[17], zll_main_rotater2219_in[25], zll_main_rotater2219_in[24], zll_main_rotater2219_in[23], zll_main_rotater2219_in[22], zll_main_rotater2219_in[21], zll_main_rotater2219_in[20], zll_main_rotater2219_in[19], zll_main_rotater2219_in[18], zll_main_rotater2219_in[16], zll_main_rotater2219_in[15], zll_main_rotater2219_in[14], zll_main_rotater2219_in[13], zll_main_rotater2219_in[12], zll_main_rotater2219_in[11], zll_main_rotater2219_in[10], zll_main_rotater2219_in[9], zll_main_rotater2219_in[8], zll_main_rotater2219_in[7], zll_main_rotater2219_in[6], zll_main_rotater2219_in[5], zll_main_rotater2219_in[4], zll_main_rotater2219_in[3], zll_main_rotater2219_in[2], zll_main_rotater2219_in[1], zll_main_rotater2219_in[0]};
  assign zll_main_rotater229_in = {zll_main_rotater2222_in[31], zll_main_rotater2222_in[30], zll_main_rotater2222_in[29], zll_main_rotater2222_in[28], zll_main_rotater2222_in[27], zll_main_rotater2222_in[26], zll_main_rotater2222_in[25], zll_main_rotater2222_in[16], zll_main_rotater2222_in[24], zll_main_rotater2222_in[23], zll_main_rotater2222_in[22], zll_main_rotater2222_in[21], zll_main_rotater2222_in[20], zll_main_rotater2222_in[19], zll_main_rotater2222_in[18], zll_main_rotater2222_in[17], zll_main_rotater2222_in[15], zll_main_rotater2222_in[14], zll_main_rotater2222_in[13], zll_main_rotater2222_in[12], zll_main_rotater2222_in[11], zll_main_rotater2222_in[10], zll_main_rotater2222_in[9], zll_main_rotater2222_in[8], zll_main_rotater2222_in[7], zll_main_rotater2222_in[6], zll_main_rotater2222_in[5], zll_main_rotater2222_in[4], zll_main_rotater2222_in[3], zll_main_rotater2222_in[2], zll_main_rotater2222_in[1], zll_main_rotater2222_in[0]};
  assign zll_main_rotater228_in = {zll_main_rotater229_in[31], zll_main_rotater229_in[30], zll_main_rotater229_in[29], zll_main_rotater229_in[28], zll_main_rotater229_in[27], zll_main_rotater229_in[26], zll_main_rotater229_in[25], zll_main_rotater229_in[24], zll_main_rotater229_in[23], zll_main_rotater229_in[22], zll_main_rotater229_in[21], zll_main_rotater229_in[20], zll_main_rotater229_in[19], zll_main_rotater229_in[15], zll_main_rotater229_in[18], zll_main_rotater229_in[17], zll_main_rotater229_in[16], zll_main_rotater229_in[14], zll_main_rotater229_in[13], zll_main_rotater229_in[12], zll_main_rotater229_in[11], zll_main_rotater229_in[10], zll_main_rotater229_in[9], zll_main_rotater229_in[8], zll_main_rotater229_in[7], zll_main_rotater229_in[6], zll_main_rotater229_in[5], zll_main_rotater229_in[4], zll_main_rotater229_in[3], zll_main_rotater229_in[2], zll_main_rotater229_in[1], zll_main_rotater229_in[0]};
  assign zll_main_rotater22_in = {zll_main_rotater228_in[31], zll_main_rotater228_in[30], zll_main_rotater228_in[29], zll_main_rotater228_in[28], zll_main_rotater228_in[27], zll_main_rotater228_in[26], zll_main_rotater228_in[25], zll_main_rotater228_in[24], zll_main_rotater228_in[23], zll_main_rotater228_in[14], zll_main_rotater228_in[22], zll_main_rotater228_in[21], zll_main_rotater228_in[20], zll_main_rotater228_in[19], zll_main_rotater228_in[18], zll_main_rotater228_in[17], zll_main_rotater228_in[16], zll_main_rotater228_in[15], zll_main_rotater228_in[13], zll_main_rotater228_in[12], zll_main_rotater228_in[11], zll_main_rotater228_in[10], zll_main_rotater228_in[9], zll_main_rotater228_in[8], zll_main_rotater228_in[7], zll_main_rotater228_in[6], zll_main_rotater228_in[5], zll_main_rotater228_in[4], zll_main_rotater228_in[3], zll_main_rotater228_in[2], zll_main_rotater228_in[1], zll_main_rotater228_in[0]};
  assign zll_main_rotater223_in = {zll_main_rotater22_in[31], zll_main_rotater22_in[30], zll_main_rotater22_in[29], zll_main_rotater22_in[28], zll_main_rotater22_in[27], zll_main_rotater22_in[26], zll_main_rotater22_in[25], zll_main_rotater22_in[24], zll_main_rotater22_in[23], zll_main_rotater22_in[13], zll_main_rotater22_in[22], zll_main_rotater22_in[21], zll_main_rotater22_in[20], zll_main_rotater22_in[19], zll_main_rotater22_in[18], zll_main_rotater22_in[17], zll_main_rotater22_in[16], zll_main_rotater22_in[15], zll_main_rotater22_in[14], zll_main_rotater22_in[12], zll_main_rotater22_in[11], zll_main_rotater22_in[10], zll_main_rotater22_in[9], zll_main_rotater22_in[8], zll_main_rotater22_in[7], zll_main_rotater22_in[6], zll_main_rotater22_in[5], zll_main_rotater22_in[4], zll_main_rotater22_in[3], zll_main_rotater22_in[2], zll_main_rotater22_in[1], zll_main_rotater22_in[0]};
  assign zll_main_rotater2212_in = {zll_main_rotater223_in[31], zll_main_rotater223_in[30], zll_main_rotater223_in[29], zll_main_rotater223_in[28], zll_main_rotater223_in[27], zll_main_rotater223_in[26], zll_main_rotater223_in[25], zll_main_rotater223_in[24], zll_main_rotater223_in[23], zll_main_rotater223_in[22], zll_main_rotater223_in[21], zll_main_rotater223_in[20], zll_main_rotater223_in[19], zll_main_rotater223_in[18], zll_main_rotater223_in[17], zll_main_rotater223_in[16], zll_main_rotater223_in[15], zll_main_rotater223_in[11], zll_main_rotater223_in[14], zll_main_rotater223_in[13], zll_main_rotater223_in[12], zll_main_rotater223_in[10], zll_main_rotater223_in[9], zll_main_rotater223_in[8], zll_main_rotater223_in[7], zll_main_rotater223_in[6], zll_main_rotater223_in[5], zll_main_rotater223_in[4], zll_main_rotater223_in[3], zll_main_rotater223_in[2], zll_main_rotater223_in[1], zll_main_rotater223_in[0]};
  assign zll_main_rotater2231_in = {zll_main_rotater2212_in[31], zll_main_rotater2212_in[30], zll_main_rotater2212_in[29], zll_main_rotater2212_in[28], zll_main_rotater2212_in[27], zll_main_rotater2212_in[26], zll_main_rotater2212_in[25], zll_main_rotater2212_in[10], zll_main_rotater2212_in[24], zll_main_rotater2212_in[23], zll_main_rotater2212_in[22], zll_main_rotater2212_in[21], zll_main_rotater2212_in[20], zll_main_rotater2212_in[19], zll_main_rotater2212_in[18], zll_main_rotater2212_in[17], zll_main_rotater2212_in[16], zll_main_rotater2212_in[15], zll_main_rotater2212_in[14], zll_main_rotater2212_in[13], zll_main_rotater2212_in[12], zll_main_rotater2212_in[11], zll_main_rotater2212_in[9], zll_main_rotater2212_in[8], zll_main_rotater2212_in[7], zll_main_rotater2212_in[6], zll_main_rotater2212_in[5], zll_main_rotater2212_in[4], zll_main_rotater2212_in[3], zll_main_rotater2212_in[2], zll_main_rotater2212_in[1], zll_main_rotater2212_in[0]};
  assign zll_main_rotater222_in = {zll_main_rotater2231_in[31], zll_main_rotater2231_in[30], zll_main_rotater2231_in[29], zll_main_rotater2231_in[28], zll_main_rotater2231_in[27], zll_main_rotater2231_in[26], zll_main_rotater2231_in[25], zll_main_rotater2231_in[24], zll_main_rotater2231_in[23], zll_main_rotater2231_in[9], zll_main_rotater2231_in[22], zll_main_rotater2231_in[21], zll_main_rotater2231_in[20], zll_main_rotater2231_in[19], zll_main_rotater2231_in[18], zll_main_rotater2231_in[17], zll_main_rotater2231_in[16], zll_main_rotater2231_in[15], zll_main_rotater2231_in[14], zll_main_rotater2231_in[13], zll_main_rotater2231_in[12], zll_main_rotater2231_in[11], zll_main_rotater2231_in[10], zll_main_rotater2231_in[8], zll_main_rotater2231_in[7], zll_main_rotater2231_in[6], zll_main_rotater2231_in[5], zll_main_rotater2231_in[4], zll_main_rotater2231_in[3], zll_main_rotater2231_in[2], zll_main_rotater2231_in[1], zll_main_rotater2231_in[0]};
  assign zll_main_rotater2227_in = {zll_main_rotater222_in[8], zll_main_rotater222_in[31], zll_main_rotater222_in[30], zll_main_rotater222_in[29], zll_main_rotater222_in[28], zll_main_rotater222_in[27], zll_main_rotater222_in[26], zll_main_rotater222_in[25], zll_main_rotater222_in[24], zll_main_rotater222_in[23], zll_main_rotater222_in[22], zll_main_rotater222_in[21], zll_main_rotater222_in[20], zll_main_rotater222_in[19], zll_main_rotater222_in[18], zll_main_rotater222_in[17], zll_main_rotater222_in[16], zll_main_rotater222_in[15], zll_main_rotater222_in[14], zll_main_rotater222_in[13], zll_main_rotater222_in[12], zll_main_rotater222_in[11], zll_main_rotater222_in[10], zll_main_rotater222_in[9], zll_main_rotater222_in[7], zll_main_rotater222_in[6], zll_main_rotater222_in[5], zll_main_rotater222_in[4], zll_main_rotater222_in[3], zll_main_rotater222_in[2], zll_main_rotater222_in[1], zll_main_rotater222_in[0]};
  assign zll_main_rotater2210_in = {zll_main_rotater2227_in[31], zll_main_rotater2227_in[30], zll_main_rotater2227_in[7], zll_main_rotater2227_in[29], zll_main_rotater2227_in[28], zll_main_rotater2227_in[27], zll_main_rotater2227_in[26], zll_main_rotater2227_in[25], zll_main_rotater2227_in[24], zll_main_rotater2227_in[23], zll_main_rotater2227_in[22], zll_main_rotater2227_in[21], zll_main_rotater2227_in[20], zll_main_rotater2227_in[19], zll_main_rotater2227_in[18], zll_main_rotater2227_in[17], zll_main_rotater2227_in[16], zll_main_rotater2227_in[15], zll_main_rotater2227_in[14], zll_main_rotater2227_in[13], zll_main_rotater2227_in[12], zll_main_rotater2227_in[11], zll_main_rotater2227_in[10], zll_main_rotater2227_in[9], zll_main_rotater2227_in[8], zll_main_rotater2227_in[6], zll_main_rotater2227_in[5], zll_main_rotater2227_in[4], zll_main_rotater2227_in[3], zll_main_rotater2227_in[2], zll_main_rotater2227_in[1], zll_main_rotater2227_in[0]};
  assign zll_main_rotater225_in = {zll_main_rotater2210_in[31], zll_main_rotater2210_in[6], zll_main_rotater2210_in[30], zll_main_rotater2210_in[29], zll_main_rotater2210_in[28], zll_main_rotater2210_in[27], zll_main_rotater2210_in[26], zll_main_rotater2210_in[25], zll_main_rotater2210_in[24], zll_main_rotater2210_in[23], zll_main_rotater2210_in[22], zll_main_rotater2210_in[21], zll_main_rotater2210_in[20], zll_main_rotater2210_in[19], zll_main_rotater2210_in[18], zll_main_rotater2210_in[17], zll_main_rotater2210_in[16], zll_main_rotater2210_in[15], zll_main_rotater2210_in[14], zll_main_rotater2210_in[13], zll_main_rotater2210_in[12], zll_main_rotater2210_in[11], zll_main_rotater2210_in[10], zll_main_rotater2210_in[9], zll_main_rotater2210_in[8], zll_main_rotater2210_in[7], zll_main_rotater2210_in[5], zll_main_rotater2210_in[4], zll_main_rotater2210_in[3], zll_main_rotater2210_in[2], zll_main_rotater2210_in[1], zll_main_rotater2210_in[0]};
  assign zll_main_rotater226_in = {zll_main_rotater225_in[31], zll_main_rotater225_in[30], zll_main_rotater225_in[29], zll_main_rotater225_in[28], zll_main_rotater225_in[27], zll_main_rotater225_in[26], zll_main_rotater225_in[25], zll_main_rotater225_in[24], zll_main_rotater225_in[23], zll_main_rotater225_in[22], zll_main_rotater225_in[21], zll_main_rotater225_in[20], zll_main_rotater225_in[19], zll_main_rotater225_in[18], zll_main_rotater225_in[17], zll_main_rotater225_in[16], zll_main_rotater225_in[15], zll_main_rotater225_in[14], zll_main_rotater225_in[13], zll_main_rotater225_in[12], zll_main_rotater225_in[11], zll_main_rotater225_in[10], zll_main_rotater225_in[5], zll_main_rotater225_in[9], zll_main_rotater225_in[8], zll_main_rotater225_in[7], zll_main_rotater225_in[6], zll_main_rotater225_in[4], zll_main_rotater225_in[3], zll_main_rotater225_in[2], zll_main_rotater225_in[1], zll_main_rotater225_in[0]};
  assign zll_main_rotater2216_in = {zll_main_rotater226_in[31], zll_main_rotater226_in[30], zll_main_rotater226_in[29], zll_main_rotater226_in[28], zll_main_rotater226_in[27], zll_main_rotater226_in[26], zll_main_rotater226_in[4], zll_main_rotater226_in[25], zll_main_rotater226_in[24], zll_main_rotater226_in[23], zll_main_rotater226_in[22], zll_main_rotater226_in[21], zll_main_rotater226_in[20], zll_main_rotater226_in[19], zll_main_rotater226_in[18], zll_main_rotater226_in[17], zll_main_rotater226_in[16], zll_main_rotater226_in[15], zll_main_rotater226_in[14], zll_main_rotater226_in[13], zll_main_rotater226_in[12], zll_main_rotater226_in[11], zll_main_rotater226_in[10], zll_main_rotater226_in[9], zll_main_rotater226_in[8], zll_main_rotater226_in[7], zll_main_rotater226_in[6], zll_main_rotater226_in[5], zll_main_rotater226_in[3], zll_main_rotater226_in[2], zll_main_rotater226_in[1], zll_main_rotater226_in[0]};
  assign zll_main_rotater2220_in = {zll_main_rotater2216_in[31], zll_main_rotater2216_in[30], zll_main_rotater2216_in[29], zll_main_rotater2216_in[28], zll_main_rotater2216_in[27], zll_main_rotater2216_in[26], zll_main_rotater2216_in[25], zll_main_rotater2216_in[24], zll_main_rotater2216_in[23], zll_main_rotater2216_in[22], zll_main_rotater2216_in[21], zll_main_rotater2216_in[20], zll_main_rotater2216_in[19], zll_main_rotater2216_in[18], zll_main_rotater2216_in[17], zll_main_rotater2216_in[16], zll_main_rotater2216_in[15], zll_main_rotater2216_in[14], zll_main_rotater2216_in[13], zll_main_rotater2216_in[3], zll_main_rotater2216_in[12], zll_main_rotater2216_in[11], zll_main_rotater2216_in[10], zll_main_rotater2216_in[9], zll_main_rotater2216_in[8], zll_main_rotater2216_in[7], zll_main_rotater2216_in[6], zll_main_rotater2216_in[5], zll_main_rotater2216_in[4], zll_main_rotater2216_in[2], zll_main_rotater2216_in[1], zll_main_rotater2216_in[0]};
  assign zll_main_rotater2217_in = {zll_main_rotater2220_in[31], zll_main_rotater2220_in[30], zll_main_rotater2220_in[29], zll_main_rotater2220_in[28], zll_main_rotater2220_in[2], zll_main_rotater2220_in[27], zll_main_rotater2220_in[26], zll_main_rotater2220_in[25], zll_main_rotater2220_in[24], zll_main_rotater2220_in[23], zll_main_rotater2220_in[22], zll_main_rotater2220_in[21], zll_main_rotater2220_in[20], zll_main_rotater2220_in[19], zll_main_rotater2220_in[18], zll_main_rotater2220_in[17], zll_main_rotater2220_in[16], zll_main_rotater2220_in[15], zll_main_rotater2220_in[14], zll_main_rotater2220_in[13], zll_main_rotater2220_in[12], zll_main_rotater2220_in[11], zll_main_rotater2220_in[10], zll_main_rotater2220_in[9], zll_main_rotater2220_in[8], zll_main_rotater2220_in[7], zll_main_rotater2220_in[6], zll_main_rotater2220_in[5], zll_main_rotater2220_in[4], zll_main_rotater2220_in[3], zll_main_rotater2220_in[1], zll_main_rotater2220_in[0]};
  assign zll_main_rotater2221_in = {zll_main_rotater2217_in[31], zll_main_rotater2217_in[30], zll_main_rotater2217_in[29], zll_main_rotater2217_in[28], zll_main_rotater2217_in[27], zll_main_rotater2217_in[26], zll_main_rotater2217_in[25], zll_main_rotater2217_in[24], zll_main_rotater2217_in[1], zll_main_rotater2217_in[23], zll_main_rotater2217_in[22], zll_main_rotater2217_in[21], zll_main_rotater2217_in[20], zll_main_rotater2217_in[19], zll_main_rotater2217_in[18], zll_main_rotater2217_in[17], zll_main_rotater2217_in[16], zll_main_rotater2217_in[15], zll_main_rotater2217_in[14], zll_main_rotater2217_in[13], zll_main_rotater2217_in[12], zll_main_rotater2217_in[11], zll_main_rotater2217_in[10], zll_main_rotater2217_in[9], zll_main_rotater2217_in[8], zll_main_rotater2217_in[7], zll_main_rotater2217_in[6], zll_main_rotater2217_in[5], zll_main_rotater2217_in[4], zll_main_rotater2217_in[3], zll_main_rotater2217_in[2], zll_main_rotater2217_in[0]};
  assign xorw32_inR5 = {extresR11, {zll_main_rotater2221_in[21], zll_main_rotater2221_in[6], zll_main_rotater2221_in[22], zll_main_rotater2221_in[20], zll_main_rotater2221_in[19], zll_main_rotater2221_in[17], zll_main_rotater2221_in[7], zll_main_rotater2221_in[13], zll_main_rotater2221_in[14], zll_main_rotater2221_in[1], zll_main_rotater2221_in[4], zll_main_rotater2221_in[18], zll_main_rotater2221_in[16], zll_main_rotater2221_in[31], zll_main_rotater2221_in[28], zll_main_rotater2221_in[30], zll_main_rotater2221_in[5], zll_main_rotater2221_in[24], zll_main_rotater2221_in[10], zll_main_rotater2221_in[27], zll_main_rotater2221_in[23], zll_main_rotater2221_in[0], zll_main_rotater2221_in[9], zll_main_rotater2221_in[8], zll_main_rotater2221_in[25], zll_main_rotater2221_in[29], zll_main_rotater2221_in[15], zll_main_rotater2221_in[2], zll_main_rotater2221_in[12], zll_main_rotater2221_in[26], zll_main_rotater2221_in[3], zll_main_rotater2221_in[11]}};
  xorW32  instR14 (xorw32_inR5[63:32], xorw32_inR5[31:0], extresR12[31:0]);
  assign main_maj_in = {zll_main_step2566_in[287:256], zll_main_step2566_in[159:128], zll_main_step2566_in[63:32]};
  assign andw32_in = {main_maj_in[95:64], main_maj_in[63:32]};
  andW32  instR15 (andw32_in[63:32], andw32_in[31:0], extresR13[31:0]);
  assign andw32_inR1 = {main_maj_in[95:64], main_maj_in[31:0]};
  andW32  instR16 (andw32_inR1[63:32], andw32_inR1[31:0], extresR14[31:0]);
  assign xorw32_inR6 = {extresR13, extresR14};
  xorW32  instR17 (xorw32_inR6[63:32], xorw32_inR6[31:0], extresR15[31:0]);
  assign andw32_inR2 = {main_maj_in[63:32], main_maj_in[31:0]};
  andW32  instR18 (andw32_inR2[63:32], andw32_inR2[31:0], extresR16[31:0]);
  assign xorw32_inR7 = {extresR15, extresR16};
  xorW32  instR19 (xorw32_inR7[63:32], xorw32_inR7[31:0], extresR17[31:0]);
  assign plusw32_inR7 = {extresR12, extresR17};
  plusW32  instR20 (plusw32_inR7[63:32], plusw32_inR7[31:0], extresR18[31:0]);
  assign plusw32_inR8 = {extresR10, extresR18};
  plusW32  instR21 (plusw32_inR8[63:32], plusw32_inR8[31:0], extresR19[31:0]);
  assign main_bigsigma1_inR1 = zll_main_step2566_in[191:160];
  Main_bigsigma1  instR22 (main_bigsigma1_inR1[31:0], main_bigsigma1_outR1);
  assign main_ch_inR1 = {zll_main_step2566_in[191:160], zll_main_step2566_in[95:64], zll_main_step2566_in[223:192]};
  Main_ch  instR23 (main_ch_inR1[95:64], main_ch_inR1[63:32], main_ch_inR1[31:0], main_ch_outR1);
  assign plusw32_inR9 = {main_bigsigma1_outR1, main_ch_outR1};
  plusW32  instR24 (plusw32_inR9[63:32], plusw32_inR9[31:0], extresR20[31:0]);
  assign plusw32_inR10 = {zll_main_step2566_in[319:288], zll_main_step2566_in[255:224]};
  plusW32  instR25 (plusw32_inR10[63:32], plusw32_inR10[31:0], extresR21[31:0]);
  assign plusw32_inR11 = {extresR20, extresR21};
  plusW32  instR26 (plusw32_inR11[63:32], plusw32_inR11[31:0], extresR22[31:0]);
  assign plusw32_inR12 = {zll_main_step2566_in[31:0], extresR22};
  plusW32  instR27 (plusw32_inR12[63:32], plusw32_inR12[31:0], extresR23[31:0]);
  assign plusw32_inR13 = {zll_main_step2566_in[127:96], extresR23};
  plusW32  instR28 (plusw32_inR13[63:32], plusw32_inR13[31:0], extresR24[31:0]);
  assign zll_main_loop6_in = {zll_main_loop35_in[1291:1286], {extresR19, zll_main_step2566_in[287:256], zll_main_step2566_in[159:128], zll_main_step2566_in[63:32], extresR24, zll_main_step2566_in[191:160], zll_main_step2566_in[95:64], zll_main_step2566_in[223:192]}, zll_main_loop35_in[773:262], zll_main_loop35_in[261:6], zll_main_loop35_in[5:0]};
  assign zll_main_loop109_in = {zll_main_loop6_in[1035:1030], zll_main_loop6_in[1029:0]};
  assign zll_main_loop107_in = {zll_main_loop109_in[1035:1030], zll_main_loop109_in[773:262], zll_main_loop109_in[1029:774], zll_main_loop109_in[261:6], zll_main_loop109_in[5:0]};
  assign zll_main_loop84_in = {zll_main_loop107_in[1035:1030], zll_main_loop107_in[517:262], zll_main_loop107_in[1029:518], zll_main_loop107_in[261:6], zll_main_loop107_in[5:0]};
  assign main_incctr_in = zll_main_loop84_in[1035:1030];
  assign lit_inR63 = main_incctr_in[5:0];
  assign lit_inR64 = main_incctr_in[5:0];
  assign lit_inR65 = main_incctr_in[5:0];
  assign lit_inR66 = main_incctr_in[5:0];
  assign lit_inR67 = main_incctr_in[5:0];
  assign lit_inR68 = main_incctr_in[5:0];
  assign lit_inR69 = main_incctr_in[5:0];
  assign lit_inR70 = main_incctr_in[5:0];
  assign lit_inR71 = main_incctr_in[5:0];
  assign lit_inR72 = main_incctr_in[5:0];
  assign lit_inR73 = main_incctr_in[5:0];
  assign lit_inR74 = main_incctr_in[5:0];
  assign lit_inR75 = main_incctr_in[5:0];
  assign lit_inR76 = main_incctr_in[5:0];
  assign lit_inR77 = main_incctr_in[5:0];
  assign lit_inR78 = main_incctr_in[5:0];
  assign lit_inR79 = main_incctr_in[5:0];
  assign lit_inR80 = main_incctr_in[5:0];
  assign lit_inR81 = main_incctr_in[5:0];
  assign lit_inR82 = main_incctr_in[5:0];
  assign lit_inR83 = main_incctr_in[5:0];
  assign lit_inR84 = main_incctr_in[5:0];
  assign lit_inR85 = main_incctr_in[5:0];
  assign lit_inR86 = main_incctr_in[5:0];
  assign lit_inR87 = main_incctr_in[5:0];
  assign lit_inR88 = main_incctr_in[5:0];
  assign lit_inR89 = main_incctr_in[5:0];
  assign lit_inR90 = main_incctr_in[5:0];
  assign lit_inR91 = main_incctr_in[5:0];
  assign lit_inR92 = main_incctr_in[5:0];
  assign lit_inR93 = main_incctr_in[5:0];
  assign lit_inR94 = main_incctr_in[5:0];
  assign lit_inR95 = main_incctr_in[5:0];
  assign lit_inR96 = main_incctr_in[5:0];
  assign lit_inR97 = main_incctr_in[5:0];
  assign lit_inR98 = main_incctr_in[5:0];
  assign lit_inR99 = main_incctr_in[5:0];
  assign lit_inR100 = main_incctr_in[5:0];
  assign lit_inR101 = main_incctr_in[5:0];
  assign lit_inR102 = main_incctr_in[5:0];
  assign lit_inR103 = main_incctr_in[5:0];
  assign lit_inR104 = main_incctr_in[5:0];
  assign lit_inR105 = main_incctr_in[5:0];
  assign lit_inR106 = main_incctr_in[5:0];
  assign lit_inR107 = main_incctr_in[5:0];
  assign lit_inR108 = main_incctr_in[5:0];
  assign lit_inR109 = main_incctr_in[5:0];
  assign lit_inR110 = main_incctr_in[5:0];
  assign lit_inR111 = main_incctr_in[5:0];
  assign lit_inR112 = main_incctr_in[5:0];
  assign lit_inR113 = main_incctr_in[5:0];
  assign lit_inR114 = main_incctr_in[5:0];
  assign lit_inR115 = main_incctr_in[5:0];
  assign lit_inR116 = main_incctr_in[5:0];
  assign lit_inR117 = main_incctr_in[5:0];
  assign lit_inR118 = main_incctr_in[5:0];
  assign lit_inR119 = main_incctr_in[5:0];
  assign lit_inR120 = main_incctr_in[5:0];
  assign lit_inR121 = main_incctr_in[5:0];
  assign lit_inR122 = main_incctr_in[5:0];
  assign lit_inR123 = main_incctr_in[5:0];
  assign lit_inR124 = main_incctr_in[5:0];
  assign lit_inR125 = main_incctr_in[5:0];
  assign zll_main_loop108_in = {zll_main_loop84_in[1035:1030], zll_main_loop84_in[1029:774], zll_main_loop84_in[773:262], zll_main_loop84_in[261:6], (lit_inR125[5:0] == 6'h0) ? 6'h1 : ((lit_inR124[5:0] == 6'h1) ? 6'h2 : ((lit_inR123[5:0] == 6'h2) ? 6'h3 : ((lit_inR122[5:0] == 6'h3) ? 6'h4 : ((lit_inR121[5:0] == 6'h4) ? 6'h5 : ((lit_inR120[5:0] == 6'h5) ? 6'h6 : ((lit_inR119[5:0] == 6'h6) ? 6'h7 : ((lit_inR118[5:0] == 6'h7) ? 6'h8 : ((lit_inR117[5:0] == 6'h8) ? 6'h9 : ((lit_inR116[5:0] == 6'h9) ? 6'ha : ((lit_inR115[5:0] == 6'ha) ? 6'hb : ((lit_inR114[5:0] == 6'hb) ? 6'hc : ((lit_inR113[5:0] == 6'hc) ? 6'hd : ((lit_inR112[5:0] == 6'hd) ? 6'he : ((lit_inR111[5:0] == 6'he) ? 6'hf : ((lit_inR110[5:0] == 6'hf) ? 6'h10 : ((lit_inR109[5:0] == 6'h10) ? 6'h11 : ((lit_inR108[5:0] == 6'h11) ? 6'h12 : ((lit_inR107[5:0] == 6'h12) ? 6'h13 : ((lit_inR106[5:0] == 6'h13) ? 6'h14 : ((lit_inR105[5:0] == 6'h14) ? 6'h15 : ((lit_inR104[5:0] == 6'h15) ? 6'h16 : ((lit_inR103[5:0] == 6'h16) ? 6'h17 : ((lit_inR102[5:0] == 6'h17) ? 6'h18 : ((lit_inR101[5:0] == 6'h18) ? 6'h19 : ((lit_inR100[5:0] == 6'h19) ? 6'h1a : ((lit_inR99[5:0] == 6'h1a) ? 6'h1b : ((lit_inR98[5:0] == 6'h1b) ? 6'h1c : ((lit_inR97[5:0] == 6'h1c) ? 6'h1d : ((lit_inR96[5:0] == 6'h1d) ? 6'h1e : ((lit_inR95[5:0] == 6'h1e) ? 6'h1f : ((lit_inR94[5:0] == 6'h1f) ? 6'h20 : ((lit_inR93[5:0] == 6'h20) ? 6'h21 : ((lit_inR92[5:0] == 6'h21) ? 6'h22 : ((lit_inR91[5:0] == 6'h22) ? 6'h23 : ((lit_inR90[5:0] == 6'h23) ? 6'h24 : ((lit_inR89[5:0] == 6'h24) ? 6'h25 : ((lit_inR88[5:0] == 6'h25) ? 6'h26 : ((lit_inR87[5:0] == 6'h26) ? 6'h27 : ((lit_inR86[5:0] == 6'h27) ? 6'h28 : ((lit_inR85[5:0] == 6'h28) ? 6'h29 : ((lit_inR84[5:0] == 6'h29) ? 6'h2a : ((lit_inR83[5:0] == 6'h2a) ? 6'h2b : ((lit_inR82[5:0] == 6'h2b) ? 6'h2c : ((lit_inR81[5:0] == 6'h2c) ? 6'h2d : ((lit_inR80[5:0] == 6'h2d) ? 6'h2e : ((lit_inR79[5:0] == 6'h2e) ? 6'h2f : ((lit_inR78[5:0] == 6'h2f) ? 6'h30 : ((lit_inR77[5:0] == 6'h30) ? 6'h31 : ((lit_inR76[5:0] == 6'h31) ? 6'h32 : ((lit_inR75[5:0] == 6'h32) ? 6'h33 : ((lit_inR74[5:0] == 6'h33) ? 6'h34 : ((lit_inR73[5:0] == 6'h34) ? 6'h35 : ((lit_inR72[5:0] == 6'h35) ? 6'h36 : ((lit_inR71[5:0] == 6'h36) ? 6'h37 : ((lit_inR70[5:0] == 6'h37) ? 6'h38 : ((lit_inR69[5:0] == 6'h38) ? 6'h39 : ((lit_inR68[5:0] == 6'h39) ? 6'h3a : ((lit_inR67[5:0] == 6'h3a) ? 6'h3b : ((lit_inR66[5:0] == 6'h3b) ? 6'h3c : ((lit_inR65[5:0] == 6'h3c) ? 6'h3d : ((lit_inR64[5:0] == 6'h3d) ? 6'h3e : ((lit_inR63[5:0] == 6'h3e) ? 6'h3f : 6'h0))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))};
  assign zll_main_loop8_in = {zll_main_loop108_in[1035:1030], zll_main_loop108_in[1029:0]};
  assign zll_main_loop67_in = {zll_main_loop8_in[1029:774], zll_main_loop8_in[1035:1030], zll_main_loop8_in[773:262], zll_main_loop8_in[261:6], zll_main_loop8_in[5:0]};
  assign zll_main_loop55_in = {zll_main_loop67_in[773:262], zll_main_loop67_in[1035:780], zll_main_loop67_in[779:774], zll_main_loop67_in[261:6], zll_main_loop67_in[5:0]};
  assign zll_main_loop29_in = {zll_main_loop55_in[267:262], zll_main_loop55_in[523:268], zll_main_loop55_in[1035:524], zll_main_loop55_in[261:6], zll_main_loop55_in[5:0]};
  assign zll_main_loop112_in = zll_main_loop29_in[1035:0];
  assign zll_main_loop18_in = {zll_main_loop112_in[1029:774], zll_main_loop112_in[1035:1030], zll_main_loop112_in[773:262], zll_main_loop112_in[261:6], zll_main_loop112_in[5:0]};
  assign zll_main_loop122_in = {zll_main_loop18_in[773:262], zll_main_loop18_in[1035:780], zll_main_loop18_in[779:774], zll_main_loop18_in[261:6], zll_main_loop18_in[5:0]};
  assign zll_main_loop41_in = {{11'h1, {8'hfa{1'h0}}}, zll_main_loop122_in[267:262], zll_main_loop122_in[523:268], zll_main_loop122_in[1035:524], zll_main_loop122_in[261:6], zll_main_loop122_in[5:0]};
  assign zll_main_loop162_in = zll_main_loop41_in[1296:0];
  assign zll_main_loop154_in = {zll_main_loop162_in[1035:1030], zll_main_loop162_in[1029:774], zll_main_loop162_in[773:262], zll_main_loop162_in[261:6], zll_main_loop162_in[5:0]};
  assign zll_main_loop111_in = {zll_main_loop154_in[1029:774], zll_main_loop154_in[1035:1030], zll_main_loop154_in[773:262], zll_main_loop154_in[261:6], zll_main_loop154_in[5:0]};
  assign zll_main_loop79_in = {zll_main_loop111_in[779:774], zll_main_loop111_in[1035:780], zll_main_loop111_in[773:262], zll_main_loop111_in[261:6], zll_main_loop111_in[5:0]};
  assign res = {261'h180000000000000000000000000000000000000000000000000000000000000001, zll_main_loop79_in[1035:1030], zll_main_loop79_in[1029:774], zll_main_loop79_in[773:262], zll_main_loop79_in[261:6], zll_main_loop79_in[5:0]};
endmodule

module Main_bigsigma1 (input logic [31:0] arg0,
  output logic [31:0] res);
  logic [31:0] main_rotater6_in;
  logic [31:0] zll_main_rotater69_in;
  logic [31:0] zll_main_rotater62_in;
  logic [31:0] zll_main_rotater610_in;
  logic [31:0] zll_main_rotater611_in;
  logic [31:0] zll_main_rotater622_in;
  logic [31:0] zll_main_rotater627_in;
  logic [31:0] zll_main_rotater613_in;
  logic [31:0] zll_main_rotater614_in;
  logic [31:0] zll_main_rotater66_in;
  logic [31:0] zll_main_rotater65_in;
  logic [31:0] zll_main_rotater617_in;
  logic [31:0] zll_main_rotater64_in;
  logic [31:0] zll_main_rotater623_in;
  logic [31:0] zll_main_rotater615_in;
  logic [31:0] zll_main_rotater625_in;
  logic [31:0] zll_main_rotater629_in;
  logic [31:0] zll_main_rotater624_in;
  logic [31:0] zll_main_rotater621_in;
  logic [31:0] zll_main_rotater630_in;
  logic [31:0] zll_main_rotater628_in;
  logic [31:0] zll_main_rotater616_in;
  logic [31:0] zll_main_rotater63_in;
  logic [31:0] zll_main_rotater619_in;
  logic [31:0] zll_main_rotater631_in;
  logic [31:0] zll_main_rotater620_in;
  logic [31:0] zll_main_rotater61_in;
  logic [31:0] zll_main_rotater6_in;
  logic [31:0] zll_main_rotater67_in;
  logic [31:0] zll_main_rotater626_in;
  logic [31:0] main_rotater11_in;
  logic [31:0] zll_main_rotater118_in;
  logic [31:0] zll_main_rotater114_in;
  logic [31:0] zll_main_rotater1123_in;
  logic [31:0] zll_main_rotater116_in;
  logic [31:0] zll_main_rotater1110_in;
  logic [31:0] zll_main_rotater112_in;
  logic [31:0] zll_main_rotater1119_in;
  logic [31:0] zll_main_rotater1130_in;
  logic [31:0] zll_main_rotater111_in;
  logic [31:0] zll_main_rotater1111_in;
  logic [31:0] zll_main_rotater119_in;
  logic [31:0] zll_main_rotater1125_in;
  logic [31:0] zll_main_rotater1127_in;
  logic [31:0] zll_main_rotater1113_in;
  logic [31:0] zll_main_rotater1128_in;
  logic [31:0] zll_main_rotater11_in;
  logic [31:0] zll_main_rotater1118_in;
  logic [31:0] zll_main_rotater1114_in;
  logic [31:0] zll_main_rotater117_in;
  logic [31:0] zll_main_rotater1115_in;
  logic [31:0] zll_main_rotater1116_in;
  logic [31:0] zll_main_rotater113_in;
  logic [31:0] zll_main_rotater115_in;
  logic [31:0] zll_main_rotater1112_in;
  logic [31:0] zll_main_rotater1120_in;
  logic [31:0] zll_main_rotater1131_in;
  logic [63:0] xorw32_in;
  logic [31:0] extres;
  logic [31:0] main_rotater25_in;
  logic [31:0] zll_main_rotater2521_in;
  logic [31:0] zll_main_rotater2515_in;
  logic [31:0] zll_main_rotater2518_in;
  logic [31:0] zll_main_rotater2516_in;
  logic [31:0] zll_main_rotater251_in;
  logic [31:0] zll_main_rotater2526_in;
  logic [31:0] zll_main_rotater255_in;
  logic [31:0] zll_main_rotater2528_in;
  logic [31:0] zll_main_rotater2511_in;
  logic [31:0] zll_main_rotater259_in;
  logic [31:0] zll_main_rotater2510_in;
  logic [31:0] zll_main_rotater2527_in;
  logic [31:0] zll_main_rotater2525_in;
  logic [31:0] zll_main_rotater2520_in;
  logic [31:0] zll_main_rotater2512_in;
  logic [31:0] zll_main_rotater258_in;
  logic [31:0] zll_main_rotater254_in;
  logic [31:0] zll_main_rotater256_in;
  logic [31:0] zll_main_rotater253_in;
  logic [31:0] zll_main_rotater2529_in;
  logic [31:0] zll_main_rotater2519_in;
  logic [31:0] zll_main_rotater2514_in;
  logic [31:0] zll_main_rotater2531_in;
  logic [31:0] zll_main_rotater2517_in;
  logic [31:0] zll_main_rotater2522_in;
  logic [31:0] zll_main_rotater25_in;
  logic [31:0] zll_main_rotater252_in;
  logic [63:0] xorw32_inR1;
  logic [31:0] extresR1;
  assign main_rotater6_in = arg0;
  assign zll_main_rotater69_in = main_rotater6_in[31:0];
  assign zll_main_rotater62_in = {zll_main_rotater69_in[30], zll_main_rotater69_in[31], zll_main_rotater69_in[29], zll_main_rotater69_in[28], zll_main_rotater69_in[27], zll_main_rotater69_in[26], zll_main_rotater69_in[25], zll_main_rotater69_in[24], zll_main_rotater69_in[23], zll_main_rotater69_in[22], zll_main_rotater69_in[21], zll_main_rotater69_in[20], zll_main_rotater69_in[19], zll_main_rotater69_in[18], zll_main_rotater69_in[17], zll_main_rotater69_in[16], zll_main_rotater69_in[15], zll_main_rotater69_in[14], zll_main_rotater69_in[13], zll_main_rotater69_in[12], zll_main_rotater69_in[11], zll_main_rotater69_in[10], zll_main_rotater69_in[9], zll_main_rotater69_in[8], zll_main_rotater69_in[7], zll_main_rotater69_in[6], zll_main_rotater69_in[5], zll_main_rotater69_in[4], zll_main_rotater69_in[3], zll_main_rotater69_in[2], zll_main_rotater69_in[1], zll_main_rotater69_in[0]};
  assign zll_main_rotater610_in = {zll_main_rotater62_in[29], zll_main_rotater62_in[31], zll_main_rotater62_in[30], zll_main_rotater62_in[28], zll_main_rotater62_in[27], zll_main_rotater62_in[26], zll_main_rotater62_in[25], zll_main_rotater62_in[24], zll_main_rotater62_in[23], zll_main_rotater62_in[22], zll_main_rotater62_in[21], zll_main_rotater62_in[20], zll_main_rotater62_in[19], zll_main_rotater62_in[18], zll_main_rotater62_in[17], zll_main_rotater62_in[16], zll_main_rotater62_in[15], zll_main_rotater62_in[14], zll_main_rotater62_in[13], zll_main_rotater62_in[12], zll_main_rotater62_in[11], zll_main_rotater62_in[10], zll_main_rotater62_in[9], zll_main_rotater62_in[8], zll_main_rotater62_in[7], zll_main_rotater62_in[6], zll_main_rotater62_in[5], zll_main_rotater62_in[4], zll_main_rotater62_in[3], zll_main_rotater62_in[2], zll_main_rotater62_in[1], zll_main_rotater62_in[0]};
  assign zll_main_rotater611_in = {zll_main_rotater610_in[27], zll_main_rotater610_in[31], zll_main_rotater610_in[30], zll_main_rotater610_in[29], zll_main_rotater610_in[28], zll_main_rotater610_in[26], zll_main_rotater610_in[25], zll_main_rotater610_in[24], zll_main_rotater610_in[23], zll_main_rotater610_in[22], zll_main_rotater610_in[21], zll_main_rotater610_in[20], zll_main_rotater610_in[19], zll_main_rotater610_in[18], zll_main_rotater610_in[17], zll_main_rotater610_in[16], zll_main_rotater610_in[15], zll_main_rotater610_in[14], zll_main_rotater610_in[13], zll_main_rotater610_in[12], zll_main_rotater610_in[11], zll_main_rotater610_in[10], zll_main_rotater610_in[9], zll_main_rotater610_in[8], zll_main_rotater610_in[7], zll_main_rotater610_in[6], zll_main_rotater610_in[5], zll_main_rotater610_in[4], zll_main_rotater610_in[3], zll_main_rotater610_in[2], zll_main_rotater610_in[1], zll_main_rotater610_in[0]};
  assign zll_main_rotater622_in = {zll_main_rotater611_in[26], zll_main_rotater611_in[31], zll_main_rotater611_in[30], zll_main_rotater611_in[29], zll_main_rotater611_in[28], zll_main_rotater611_in[27], zll_main_rotater611_in[25], zll_main_rotater611_in[24], zll_main_rotater611_in[23], zll_main_rotater611_in[22], zll_main_rotater611_in[21], zll_main_rotater611_in[20], zll_main_rotater611_in[19], zll_main_rotater611_in[18], zll_main_rotater611_in[17], zll_main_rotater611_in[16], zll_main_rotater611_in[15], zll_main_rotater611_in[14], zll_main_rotater611_in[13], zll_main_rotater611_in[12], zll_main_rotater611_in[11], zll_main_rotater611_in[10], zll_main_rotater611_in[9], zll_main_rotater611_in[8], zll_main_rotater611_in[7], zll_main_rotater611_in[6], zll_main_rotater611_in[5], zll_main_rotater611_in[4], zll_main_rotater611_in[3], zll_main_rotater611_in[2], zll_main_rotater611_in[1], zll_main_rotater611_in[0]};
  assign zll_main_rotater627_in = {zll_main_rotater622_in[31], zll_main_rotater622_in[30], zll_main_rotater622_in[29], zll_main_rotater622_in[28], zll_main_rotater622_in[25], zll_main_rotater622_in[27], zll_main_rotater622_in[26], zll_main_rotater622_in[24], zll_main_rotater622_in[23], zll_main_rotater622_in[22], zll_main_rotater622_in[21], zll_main_rotater622_in[20], zll_main_rotater622_in[19], zll_main_rotater622_in[18], zll_main_rotater622_in[17], zll_main_rotater622_in[16], zll_main_rotater622_in[15], zll_main_rotater622_in[14], zll_main_rotater622_in[13], zll_main_rotater622_in[12], zll_main_rotater622_in[11], zll_main_rotater622_in[10], zll_main_rotater622_in[9], zll_main_rotater622_in[8], zll_main_rotater622_in[7], zll_main_rotater622_in[6], zll_main_rotater622_in[5], zll_main_rotater622_in[4], zll_main_rotater622_in[3], zll_main_rotater622_in[2], zll_main_rotater622_in[1], zll_main_rotater622_in[0]};
  assign zll_main_rotater613_in = {zll_main_rotater627_in[31], zll_main_rotater627_in[30], zll_main_rotater627_in[29], zll_main_rotater627_in[28], zll_main_rotater627_in[24], zll_main_rotater627_in[27], zll_main_rotater627_in[26], zll_main_rotater627_in[25], zll_main_rotater627_in[23], zll_main_rotater627_in[22], zll_main_rotater627_in[21], zll_main_rotater627_in[20], zll_main_rotater627_in[19], zll_main_rotater627_in[18], zll_main_rotater627_in[17], zll_main_rotater627_in[16], zll_main_rotater627_in[15], zll_main_rotater627_in[14], zll_main_rotater627_in[13], zll_main_rotater627_in[12], zll_main_rotater627_in[11], zll_main_rotater627_in[10], zll_main_rotater627_in[9], zll_main_rotater627_in[8], zll_main_rotater627_in[7], zll_main_rotater627_in[6], zll_main_rotater627_in[5], zll_main_rotater627_in[4], zll_main_rotater627_in[3], zll_main_rotater627_in[2], zll_main_rotater627_in[1], zll_main_rotater627_in[0]};
  assign zll_main_rotater614_in = {zll_main_rotater613_in[31], zll_main_rotater613_in[30], zll_main_rotater613_in[29], zll_main_rotater613_in[28], zll_main_rotater613_in[27], zll_main_rotater613_in[23], zll_main_rotater613_in[26], zll_main_rotater613_in[25], zll_main_rotater613_in[24], zll_main_rotater613_in[22], zll_main_rotater613_in[21], zll_main_rotater613_in[20], zll_main_rotater613_in[19], zll_main_rotater613_in[18], zll_main_rotater613_in[17], zll_main_rotater613_in[16], zll_main_rotater613_in[15], zll_main_rotater613_in[14], zll_main_rotater613_in[13], zll_main_rotater613_in[12], zll_main_rotater613_in[11], zll_main_rotater613_in[10], zll_main_rotater613_in[9], zll_main_rotater613_in[8], zll_main_rotater613_in[7], zll_main_rotater613_in[6], zll_main_rotater613_in[5], zll_main_rotater613_in[4], zll_main_rotater613_in[3], zll_main_rotater613_in[2], zll_main_rotater613_in[1], zll_main_rotater613_in[0]};
  assign zll_main_rotater66_in = {zll_main_rotater614_in[31], zll_main_rotater614_in[30], zll_main_rotater614_in[29], zll_main_rotater614_in[28], zll_main_rotater614_in[27], zll_main_rotater614_in[22], zll_main_rotater614_in[26], zll_main_rotater614_in[25], zll_main_rotater614_in[24], zll_main_rotater614_in[23], zll_main_rotater614_in[21], zll_main_rotater614_in[20], zll_main_rotater614_in[19], zll_main_rotater614_in[18], zll_main_rotater614_in[17], zll_main_rotater614_in[16], zll_main_rotater614_in[15], zll_main_rotater614_in[14], zll_main_rotater614_in[13], zll_main_rotater614_in[12], zll_main_rotater614_in[11], zll_main_rotater614_in[10], zll_main_rotater614_in[9], zll_main_rotater614_in[8], zll_main_rotater614_in[7], zll_main_rotater614_in[6], zll_main_rotater614_in[5], zll_main_rotater614_in[4], zll_main_rotater614_in[3], zll_main_rotater614_in[2], zll_main_rotater614_in[1], zll_main_rotater614_in[0]};
  assign zll_main_rotater65_in = {zll_main_rotater66_in[31], zll_main_rotater66_in[30], zll_main_rotater66_in[29], zll_main_rotater66_in[28], zll_main_rotater66_in[21], zll_main_rotater66_in[27], zll_main_rotater66_in[26], zll_main_rotater66_in[25], zll_main_rotater66_in[24], zll_main_rotater66_in[23], zll_main_rotater66_in[22], zll_main_rotater66_in[20], zll_main_rotater66_in[19], zll_main_rotater66_in[18], zll_main_rotater66_in[17], zll_main_rotater66_in[16], zll_main_rotater66_in[15], zll_main_rotater66_in[14], zll_main_rotater66_in[13], zll_main_rotater66_in[12], zll_main_rotater66_in[11], zll_main_rotater66_in[10], zll_main_rotater66_in[9], zll_main_rotater66_in[8], zll_main_rotater66_in[7], zll_main_rotater66_in[6], zll_main_rotater66_in[5], zll_main_rotater66_in[4], zll_main_rotater66_in[3], zll_main_rotater66_in[2], zll_main_rotater66_in[1], zll_main_rotater66_in[0]};
  assign zll_main_rotater617_in = {zll_main_rotater65_in[31], zll_main_rotater65_in[30], zll_main_rotater65_in[29], zll_main_rotater65_in[28], zll_main_rotater65_in[27], zll_main_rotater65_in[26], zll_main_rotater65_in[20], zll_main_rotater65_in[25], zll_main_rotater65_in[24], zll_main_rotater65_in[23], zll_main_rotater65_in[22], zll_main_rotater65_in[21], zll_main_rotater65_in[19], zll_main_rotater65_in[18], zll_main_rotater65_in[17], zll_main_rotater65_in[16], zll_main_rotater65_in[15], zll_main_rotater65_in[14], zll_main_rotater65_in[13], zll_main_rotater65_in[12], zll_main_rotater65_in[11], zll_main_rotater65_in[10], zll_main_rotater65_in[9], zll_main_rotater65_in[8], zll_main_rotater65_in[7], zll_main_rotater65_in[6], zll_main_rotater65_in[5], zll_main_rotater65_in[4], zll_main_rotater65_in[3], zll_main_rotater65_in[2], zll_main_rotater65_in[1], zll_main_rotater65_in[0]};
  assign zll_main_rotater64_in = {zll_main_rotater617_in[31], zll_main_rotater617_in[18], zll_main_rotater617_in[30], zll_main_rotater617_in[29], zll_main_rotater617_in[28], zll_main_rotater617_in[27], zll_main_rotater617_in[26], zll_main_rotater617_in[25], zll_main_rotater617_in[24], zll_main_rotater617_in[23], zll_main_rotater617_in[22], zll_main_rotater617_in[21], zll_main_rotater617_in[20], zll_main_rotater617_in[19], zll_main_rotater617_in[17], zll_main_rotater617_in[16], zll_main_rotater617_in[15], zll_main_rotater617_in[14], zll_main_rotater617_in[13], zll_main_rotater617_in[12], zll_main_rotater617_in[11], zll_main_rotater617_in[10], zll_main_rotater617_in[9], zll_main_rotater617_in[8], zll_main_rotater617_in[7], zll_main_rotater617_in[6], zll_main_rotater617_in[5], zll_main_rotater617_in[4], zll_main_rotater617_in[3], zll_main_rotater617_in[2], zll_main_rotater617_in[1], zll_main_rotater617_in[0]};
  assign zll_main_rotater623_in = {zll_main_rotater64_in[31], zll_main_rotater64_in[30], zll_main_rotater64_in[29], zll_main_rotater64_in[17], zll_main_rotater64_in[28], zll_main_rotater64_in[27], zll_main_rotater64_in[26], zll_main_rotater64_in[25], zll_main_rotater64_in[24], zll_main_rotater64_in[23], zll_main_rotater64_in[22], zll_main_rotater64_in[21], zll_main_rotater64_in[20], zll_main_rotater64_in[19], zll_main_rotater64_in[18], zll_main_rotater64_in[16], zll_main_rotater64_in[15], zll_main_rotater64_in[14], zll_main_rotater64_in[13], zll_main_rotater64_in[12], zll_main_rotater64_in[11], zll_main_rotater64_in[10], zll_main_rotater64_in[9], zll_main_rotater64_in[8], zll_main_rotater64_in[7], zll_main_rotater64_in[6], zll_main_rotater64_in[5], zll_main_rotater64_in[4], zll_main_rotater64_in[3], zll_main_rotater64_in[2], zll_main_rotater64_in[1], zll_main_rotater64_in[0]};
  assign zll_main_rotater615_in = {zll_main_rotater623_in[31], zll_main_rotater623_in[30], zll_main_rotater623_in[29], zll_main_rotater623_in[28], zll_main_rotater623_in[27], zll_main_rotater623_in[26], zll_main_rotater623_in[25], zll_main_rotater623_in[24], zll_main_rotater623_in[23], zll_main_rotater623_in[22], zll_main_rotater623_in[16], zll_main_rotater623_in[21], zll_main_rotater623_in[20], zll_main_rotater623_in[19], zll_main_rotater623_in[18], zll_main_rotater623_in[17], zll_main_rotater623_in[15], zll_main_rotater623_in[14], zll_main_rotater623_in[13], zll_main_rotater623_in[12], zll_main_rotater623_in[11], zll_main_rotater623_in[10], zll_main_rotater623_in[9], zll_main_rotater623_in[8], zll_main_rotater623_in[7], zll_main_rotater623_in[6], zll_main_rotater623_in[5], zll_main_rotater623_in[4], zll_main_rotater623_in[3], zll_main_rotater623_in[2], zll_main_rotater623_in[1], zll_main_rotater623_in[0]};
  assign zll_main_rotater625_in = {zll_main_rotater615_in[31], zll_main_rotater615_in[15], zll_main_rotater615_in[30], zll_main_rotater615_in[29], zll_main_rotater615_in[28], zll_main_rotater615_in[27], zll_main_rotater615_in[26], zll_main_rotater615_in[25], zll_main_rotater615_in[24], zll_main_rotater615_in[23], zll_main_rotater615_in[22], zll_main_rotater615_in[21], zll_main_rotater615_in[20], zll_main_rotater615_in[19], zll_main_rotater615_in[18], zll_main_rotater615_in[17], zll_main_rotater615_in[16], zll_main_rotater615_in[14], zll_main_rotater615_in[13], zll_main_rotater615_in[12], zll_main_rotater615_in[11], zll_main_rotater615_in[10], zll_main_rotater615_in[9], zll_main_rotater615_in[8], zll_main_rotater615_in[7], zll_main_rotater615_in[6], zll_main_rotater615_in[5], zll_main_rotater615_in[4], zll_main_rotater615_in[3], zll_main_rotater615_in[2], zll_main_rotater615_in[1], zll_main_rotater615_in[0]};
  assign zll_main_rotater629_in = {zll_main_rotater625_in[31], zll_main_rotater625_in[30], zll_main_rotater625_in[29], zll_main_rotater625_in[28], zll_main_rotater625_in[27], zll_main_rotater625_in[26], zll_main_rotater625_in[25], zll_main_rotater625_in[24], zll_main_rotater625_in[23], zll_main_rotater625_in[22], zll_main_rotater625_in[14], zll_main_rotater625_in[21], zll_main_rotater625_in[20], zll_main_rotater625_in[19], zll_main_rotater625_in[18], zll_main_rotater625_in[17], zll_main_rotater625_in[16], zll_main_rotater625_in[15], zll_main_rotater625_in[13], zll_main_rotater625_in[12], zll_main_rotater625_in[11], zll_main_rotater625_in[10], zll_main_rotater625_in[9], zll_main_rotater625_in[8], zll_main_rotater625_in[7], zll_main_rotater625_in[6], zll_main_rotater625_in[5], zll_main_rotater625_in[4], zll_main_rotater625_in[3], zll_main_rotater625_in[2], zll_main_rotater625_in[1], zll_main_rotater625_in[0]};
  assign zll_main_rotater624_in = {zll_main_rotater629_in[31], zll_main_rotater629_in[30], zll_main_rotater629_in[29], zll_main_rotater629_in[28], zll_main_rotater629_in[27], zll_main_rotater629_in[26], zll_main_rotater629_in[25], zll_main_rotater629_in[24], zll_main_rotater629_in[23], zll_main_rotater629_in[13], zll_main_rotater629_in[22], zll_main_rotater629_in[21], zll_main_rotater629_in[20], zll_main_rotater629_in[19], zll_main_rotater629_in[18], zll_main_rotater629_in[17], zll_main_rotater629_in[16], zll_main_rotater629_in[15], zll_main_rotater629_in[14], zll_main_rotater629_in[12], zll_main_rotater629_in[11], zll_main_rotater629_in[10], zll_main_rotater629_in[9], zll_main_rotater629_in[8], zll_main_rotater629_in[7], zll_main_rotater629_in[6], zll_main_rotater629_in[5], zll_main_rotater629_in[4], zll_main_rotater629_in[3], zll_main_rotater629_in[2], zll_main_rotater629_in[1], zll_main_rotater629_in[0]};
  assign zll_main_rotater621_in = {zll_main_rotater624_in[31], zll_main_rotater624_in[30], zll_main_rotater624_in[29], zll_main_rotater624_in[28], zll_main_rotater624_in[27], zll_main_rotater624_in[26], zll_main_rotater624_in[25], zll_main_rotater624_in[24], zll_main_rotater624_in[23], zll_main_rotater624_in[22], zll_main_rotater624_in[21], zll_main_rotater624_in[20], zll_main_rotater624_in[19], zll_main_rotater624_in[18], zll_main_rotater624_in[17], zll_main_rotater624_in[16], zll_main_rotater624_in[12], zll_main_rotater624_in[15], zll_main_rotater624_in[14], zll_main_rotater624_in[13], zll_main_rotater624_in[11], zll_main_rotater624_in[10], zll_main_rotater624_in[9], zll_main_rotater624_in[8], zll_main_rotater624_in[7], zll_main_rotater624_in[6], zll_main_rotater624_in[5], zll_main_rotater624_in[4], zll_main_rotater624_in[3], zll_main_rotater624_in[2], zll_main_rotater624_in[1], zll_main_rotater624_in[0]};
  assign zll_main_rotater630_in = {zll_main_rotater621_in[31], zll_main_rotater621_in[30], zll_main_rotater621_in[29], zll_main_rotater621_in[28], zll_main_rotater621_in[27], zll_main_rotater621_in[11], zll_main_rotater621_in[26], zll_main_rotater621_in[25], zll_main_rotater621_in[24], zll_main_rotater621_in[23], zll_main_rotater621_in[22], zll_main_rotater621_in[21], zll_main_rotater621_in[20], zll_main_rotater621_in[19], zll_main_rotater621_in[18], zll_main_rotater621_in[17], zll_main_rotater621_in[16], zll_main_rotater621_in[15], zll_main_rotater621_in[14], zll_main_rotater621_in[13], zll_main_rotater621_in[12], zll_main_rotater621_in[10], zll_main_rotater621_in[9], zll_main_rotater621_in[8], zll_main_rotater621_in[7], zll_main_rotater621_in[6], zll_main_rotater621_in[5], zll_main_rotater621_in[4], zll_main_rotater621_in[3], zll_main_rotater621_in[2], zll_main_rotater621_in[1], zll_main_rotater621_in[0]};
  assign zll_main_rotater628_in = {zll_main_rotater630_in[10], zll_main_rotater630_in[31], zll_main_rotater630_in[30], zll_main_rotater630_in[29], zll_main_rotater630_in[28], zll_main_rotater630_in[27], zll_main_rotater630_in[26], zll_main_rotater630_in[25], zll_main_rotater630_in[24], zll_main_rotater630_in[23], zll_main_rotater630_in[22], zll_main_rotater630_in[21], zll_main_rotater630_in[20], zll_main_rotater630_in[19], zll_main_rotater630_in[18], zll_main_rotater630_in[17], zll_main_rotater630_in[16], zll_main_rotater630_in[15], zll_main_rotater630_in[14], zll_main_rotater630_in[13], zll_main_rotater630_in[12], zll_main_rotater630_in[11], zll_main_rotater630_in[9], zll_main_rotater630_in[8], zll_main_rotater630_in[7], zll_main_rotater630_in[6], zll_main_rotater630_in[5], zll_main_rotater630_in[4], zll_main_rotater630_in[3], zll_main_rotater630_in[2], zll_main_rotater630_in[1], zll_main_rotater630_in[0]};
  assign zll_main_rotater616_in = {zll_main_rotater628_in[31], zll_main_rotater628_in[9], zll_main_rotater628_in[30], zll_main_rotater628_in[29], zll_main_rotater628_in[28], zll_main_rotater628_in[27], zll_main_rotater628_in[26], zll_main_rotater628_in[25], zll_main_rotater628_in[24], zll_main_rotater628_in[23], zll_main_rotater628_in[22], zll_main_rotater628_in[21], zll_main_rotater628_in[20], zll_main_rotater628_in[19], zll_main_rotater628_in[18], zll_main_rotater628_in[17], zll_main_rotater628_in[16], zll_main_rotater628_in[15], zll_main_rotater628_in[14], zll_main_rotater628_in[13], zll_main_rotater628_in[12], zll_main_rotater628_in[11], zll_main_rotater628_in[10], zll_main_rotater628_in[8], zll_main_rotater628_in[7], zll_main_rotater628_in[6], zll_main_rotater628_in[5], zll_main_rotater628_in[4], zll_main_rotater628_in[3], zll_main_rotater628_in[2], zll_main_rotater628_in[1], zll_main_rotater628_in[0]};
  assign zll_main_rotater63_in = {zll_main_rotater616_in[31], zll_main_rotater616_in[30], zll_main_rotater616_in[29], zll_main_rotater616_in[28], zll_main_rotater616_in[27], zll_main_rotater616_in[26], zll_main_rotater616_in[25], zll_main_rotater616_in[24], zll_main_rotater616_in[23], zll_main_rotater616_in[22], zll_main_rotater616_in[21], zll_main_rotater616_in[20], zll_main_rotater616_in[19], zll_main_rotater616_in[18], zll_main_rotater616_in[17], zll_main_rotater616_in[16], zll_main_rotater616_in[15], zll_main_rotater616_in[14], zll_main_rotater616_in[13], zll_main_rotater616_in[8], zll_main_rotater616_in[12], zll_main_rotater616_in[11], zll_main_rotater616_in[10], zll_main_rotater616_in[9], zll_main_rotater616_in[7], zll_main_rotater616_in[6], zll_main_rotater616_in[5], zll_main_rotater616_in[4], zll_main_rotater616_in[3], zll_main_rotater616_in[2], zll_main_rotater616_in[1], zll_main_rotater616_in[0]};
  assign zll_main_rotater619_in = {zll_main_rotater63_in[31], zll_main_rotater63_in[30], zll_main_rotater63_in[29], zll_main_rotater63_in[7], zll_main_rotater63_in[28], zll_main_rotater63_in[27], zll_main_rotater63_in[26], zll_main_rotater63_in[25], zll_main_rotater63_in[24], zll_main_rotater63_in[23], zll_main_rotater63_in[22], zll_main_rotater63_in[21], zll_main_rotater63_in[20], zll_main_rotater63_in[19], zll_main_rotater63_in[18], zll_main_rotater63_in[17], zll_main_rotater63_in[16], zll_main_rotater63_in[15], zll_main_rotater63_in[14], zll_main_rotater63_in[13], zll_main_rotater63_in[12], zll_main_rotater63_in[11], zll_main_rotater63_in[10], zll_main_rotater63_in[9], zll_main_rotater63_in[8], zll_main_rotater63_in[6], zll_main_rotater63_in[5], zll_main_rotater63_in[4], zll_main_rotater63_in[3], zll_main_rotater63_in[2], zll_main_rotater63_in[1], zll_main_rotater63_in[0]};
  assign zll_main_rotater631_in = {zll_main_rotater619_in[31], zll_main_rotater619_in[30], zll_main_rotater619_in[6], zll_main_rotater619_in[29], zll_main_rotater619_in[28], zll_main_rotater619_in[27], zll_main_rotater619_in[26], zll_main_rotater619_in[25], zll_main_rotater619_in[24], zll_main_rotater619_in[23], zll_main_rotater619_in[22], zll_main_rotater619_in[21], zll_main_rotater619_in[20], zll_main_rotater619_in[19], zll_main_rotater619_in[18], zll_main_rotater619_in[17], zll_main_rotater619_in[16], zll_main_rotater619_in[15], zll_main_rotater619_in[14], zll_main_rotater619_in[13], zll_main_rotater619_in[12], zll_main_rotater619_in[11], zll_main_rotater619_in[10], zll_main_rotater619_in[9], zll_main_rotater619_in[8], zll_main_rotater619_in[7], zll_main_rotater619_in[5], zll_main_rotater619_in[4], zll_main_rotater619_in[3], zll_main_rotater619_in[2], zll_main_rotater619_in[1], zll_main_rotater619_in[0]};
  assign zll_main_rotater620_in = {zll_main_rotater631_in[31], zll_main_rotater631_in[30], zll_main_rotater631_in[29], zll_main_rotater631_in[5], zll_main_rotater631_in[28], zll_main_rotater631_in[27], zll_main_rotater631_in[26], zll_main_rotater631_in[25], zll_main_rotater631_in[24], zll_main_rotater631_in[23], zll_main_rotater631_in[22], zll_main_rotater631_in[21], zll_main_rotater631_in[20], zll_main_rotater631_in[19], zll_main_rotater631_in[18], zll_main_rotater631_in[17], zll_main_rotater631_in[16], zll_main_rotater631_in[15], zll_main_rotater631_in[14], zll_main_rotater631_in[13], zll_main_rotater631_in[12], zll_main_rotater631_in[11], zll_main_rotater631_in[10], zll_main_rotater631_in[9], zll_main_rotater631_in[8], zll_main_rotater631_in[7], zll_main_rotater631_in[6], zll_main_rotater631_in[4], zll_main_rotater631_in[3], zll_main_rotater631_in[2], zll_main_rotater631_in[1], zll_main_rotater631_in[0]};
  assign zll_main_rotater61_in = {zll_main_rotater620_in[31], zll_main_rotater620_in[30], zll_main_rotater620_in[29], zll_main_rotater620_in[28], zll_main_rotater620_in[27], zll_main_rotater620_in[26], zll_main_rotater620_in[25], zll_main_rotater620_in[24], zll_main_rotater620_in[4], zll_main_rotater620_in[23], zll_main_rotater620_in[22], zll_main_rotater620_in[21], zll_main_rotater620_in[20], zll_main_rotater620_in[19], zll_main_rotater620_in[18], zll_main_rotater620_in[17], zll_main_rotater620_in[16], zll_main_rotater620_in[15], zll_main_rotater620_in[14], zll_main_rotater620_in[13], zll_main_rotater620_in[12], zll_main_rotater620_in[11], zll_main_rotater620_in[10], zll_main_rotater620_in[9], zll_main_rotater620_in[8], zll_main_rotater620_in[7], zll_main_rotater620_in[6], zll_main_rotater620_in[5], zll_main_rotater620_in[3], zll_main_rotater620_in[2], zll_main_rotater620_in[1], zll_main_rotater620_in[0]};
  assign zll_main_rotater6_in = {zll_main_rotater61_in[31], zll_main_rotater61_in[30], zll_main_rotater61_in[29], zll_main_rotater61_in[28], zll_main_rotater61_in[27], zll_main_rotater61_in[26], zll_main_rotater61_in[25], zll_main_rotater61_in[24], zll_main_rotater61_in[23], zll_main_rotater61_in[22], zll_main_rotater61_in[21], zll_main_rotater61_in[20], zll_main_rotater61_in[19], zll_main_rotater61_in[18], zll_main_rotater61_in[17], zll_main_rotater61_in[16], zll_main_rotater61_in[15], zll_main_rotater61_in[14], zll_main_rotater61_in[13], zll_main_rotater61_in[12], zll_main_rotater61_in[11], zll_main_rotater61_in[10], zll_main_rotater61_in[9], zll_main_rotater61_in[8], zll_main_rotater61_in[7], zll_main_rotater61_in[3], zll_main_rotater61_in[6], zll_main_rotater61_in[5], zll_main_rotater61_in[4], zll_main_rotater61_in[2], zll_main_rotater61_in[1], zll_main_rotater61_in[0]};
  assign zll_main_rotater67_in = {zll_main_rotater6_in[31], zll_main_rotater6_in[30], zll_main_rotater6_in[29], zll_main_rotater6_in[28], zll_main_rotater6_in[27], zll_main_rotater6_in[26], zll_main_rotater6_in[2], zll_main_rotater6_in[25], zll_main_rotater6_in[24], zll_main_rotater6_in[23], zll_main_rotater6_in[22], zll_main_rotater6_in[21], zll_main_rotater6_in[20], zll_main_rotater6_in[19], zll_main_rotater6_in[18], zll_main_rotater6_in[17], zll_main_rotater6_in[16], zll_main_rotater6_in[15], zll_main_rotater6_in[14], zll_main_rotater6_in[13], zll_main_rotater6_in[12], zll_main_rotater6_in[11], zll_main_rotater6_in[10], zll_main_rotater6_in[9], zll_main_rotater6_in[8], zll_main_rotater6_in[7], zll_main_rotater6_in[6], zll_main_rotater6_in[5], zll_main_rotater6_in[4], zll_main_rotater6_in[3], zll_main_rotater6_in[1], zll_main_rotater6_in[0]};
  assign zll_main_rotater626_in = {zll_main_rotater67_in[31], zll_main_rotater67_in[30], zll_main_rotater67_in[29], zll_main_rotater67_in[28], zll_main_rotater67_in[27], zll_main_rotater67_in[26], zll_main_rotater67_in[25], zll_main_rotater67_in[24], zll_main_rotater67_in[23], zll_main_rotater67_in[22], zll_main_rotater67_in[21], zll_main_rotater67_in[20], zll_main_rotater67_in[19], zll_main_rotater67_in[18], zll_main_rotater67_in[17], zll_main_rotater67_in[1], zll_main_rotater67_in[16], zll_main_rotater67_in[15], zll_main_rotater67_in[14], zll_main_rotater67_in[13], zll_main_rotater67_in[12], zll_main_rotater67_in[11], zll_main_rotater67_in[10], zll_main_rotater67_in[9], zll_main_rotater67_in[8], zll_main_rotater67_in[7], zll_main_rotater67_in[6], zll_main_rotater67_in[5], zll_main_rotater67_in[4], zll_main_rotater67_in[3], zll_main_rotater67_in[2], zll_main_rotater67_in[0]};
  assign main_rotater11_in = arg0;
  assign zll_main_rotater118_in = main_rotater11_in[31:0];
  assign zll_main_rotater114_in = {zll_main_rotater118_in[31], zll_main_rotater118_in[29], zll_main_rotater118_in[30], zll_main_rotater118_in[28], zll_main_rotater118_in[27], zll_main_rotater118_in[26], zll_main_rotater118_in[25], zll_main_rotater118_in[24], zll_main_rotater118_in[23], zll_main_rotater118_in[22], zll_main_rotater118_in[21], zll_main_rotater118_in[20], zll_main_rotater118_in[19], zll_main_rotater118_in[18], zll_main_rotater118_in[17], zll_main_rotater118_in[16], zll_main_rotater118_in[15], zll_main_rotater118_in[14], zll_main_rotater118_in[13], zll_main_rotater118_in[12], zll_main_rotater118_in[11], zll_main_rotater118_in[10], zll_main_rotater118_in[9], zll_main_rotater118_in[8], zll_main_rotater118_in[7], zll_main_rotater118_in[6], zll_main_rotater118_in[5], zll_main_rotater118_in[4], zll_main_rotater118_in[3], zll_main_rotater118_in[2], zll_main_rotater118_in[1], zll_main_rotater118_in[0]};
  assign zll_main_rotater1123_in = {zll_main_rotater114_in[28], zll_main_rotater114_in[31], zll_main_rotater114_in[30], zll_main_rotater114_in[29], zll_main_rotater114_in[27], zll_main_rotater114_in[26], zll_main_rotater114_in[25], zll_main_rotater114_in[24], zll_main_rotater114_in[23], zll_main_rotater114_in[22], zll_main_rotater114_in[21], zll_main_rotater114_in[20], zll_main_rotater114_in[19], zll_main_rotater114_in[18], zll_main_rotater114_in[17], zll_main_rotater114_in[16], zll_main_rotater114_in[15], zll_main_rotater114_in[14], zll_main_rotater114_in[13], zll_main_rotater114_in[12], zll_main_rotater114_in[11], zll_main_rotater114_in[10], zll_main_rotater114_in[9], zll_main_rotater114_in[8], zll_main_rotater114_in[7], zll_main_rotater114_in[6], zll_main_rotater114_in[5], zll_main_rotater114_in[4], zll_main_rotater114_in[3], zll_main_rotater114_in[2], zll_main_rotater114_in[1], zll_main_rotater114_in[0]};
  assign zll_main_rotater116_in = {zll_main_rotater1123_in[31], zll_main_rotater1123_in[30], zll_main_rotater1123_in[29], zll_main_rotater1123_in[27], zll_main_rotater1123_in[28], zll_main_rotater1123_in[26], zll_main_rotater1123_in[25], zll_main_rotater1123_in[24], zll_main_rotater1123_in[23], zll_main_rotater1123_in[22], zll_main_rotater1123_in[21], zll_main_rotater1123_in[20], zll_main_rotater1123_in[19], zll_main_rotater1123_in[18], zll_main_rotater1123_in[17], zll_main_rotater1123_in[16], zll_main_rotater1123_in[15], zll_main_rotater1123_in[14], zll_main_rotater1123_in[13], zll_main_rotater1123_in[12], zll_main_rotater1123_in[11], zll_main_rotater1123_in[10], zll_main_rotater1123_in[9], zll_main_rotater1123_in[8], zll_main_rotater1123_in[7], zll_main_rotater1123_in[6], zll_main_rotater1123_in[5], zll_main_rotater1123_in[4], zll_main_rotater1123_in[3], zll_main_rotater1123_in[2], zll_main_rotater1123_in[1], zll_main_rotater1123_in[0]};
  assign zll_main_rotater1110_in = {zll_main_rotater116_in[24], zll_main_rotater116_in[31], zll_main_rotater116_in[30], zll_main_rotater116_in[29], zll_main_rotater116_in[28], zll_main_rotater116_in[27], zll_main_rotater116_in[26], zll_main_rotater116_in[25], zll_main_rotater116_in[23], zll_main_rotater116_in[22], zll_main_rotater116_in[21], zll_main_rotater116_in[20], zll_main_rotater116_in[19], zll_main_rotater116_in[18], zll_main_rotater116_in[17], zll_main_rotater116_in[16], zll_main_rotater116_in[15], zll_main_rotater116_in[14], zll_main_rotater116_in[13], zll_main_rotater116_in[12], zll_main_rotater116_in[11], zll_main_rotater116_in[10], zll_main_rotater116_in[9], zll_main_rotater116_in[8], zll_main_rotater116_in[7], zll_main_rotater116_in[6], zll_main_rotater116_in[5], zll_main_rotater116_in[4], zll_main_rotater116_in[3], zll_main_rotater116_in[2], zll_main_rotater116_in[1], zll_main_rotater116_in[0]};
  assign zll_main_rotater112_in = {zll_main_rotater1110_in[23], zll_main_rotater1110_in[31], zll_main_rotater1110_in[30], zll_main_rotater1110_in[29], zll_main_rotater1110_in[28], zll_main_rotater1110_in[27], zll_main_rotater1110_in[26], zll_main_rotater1110_in[25], zll_main_rotater1110_in[24], zll_main_rotater1110_in[22], zll_main_rotater1110_in[21], zll_main_rotater1110_in[20], zll_main_rotater1110_in[19], zll_main_rotater1110_in[18], zll_main_rotater1110_in[17], zll_main_rotater1110_in[16], zll_main_rotater1110_in[15], zll_main_rotater1110_in[14], zll_main_rotater1110_in[13], zll_main_rotater1110_in[12], zll_main_rotater1110_in[11], zll_main_rotater1110_in[10], zll_main_rotater1110_in[9], zll_main_rotater1110_in[8], zll_main_rotater1110_in[7], zll_main_rotater1110_in[6], zll_main_rotater1110_in[5], zll_main_rotater1110_in[4], zll_main_rotater1110_in[3], zll_main_rotater1110_in[2], zll_main_rotater1110_in[1], zll_main_rotater1110_in[0]};
  assign zll_main_rotater1119_in = {zll_main_rotater112_in[31], zll_main_rotater112_in[30], zll_main_rotater112_in[29], zll_main_rotater112_in[28], zll_main_rotater112_in[27], zll_main_rotater112_in[26], zll_main_rotater112_in[25], zll_main_rotater112_in[24], zll_main_rotater112_in[21], zll_main_rotater112_in[23], zll_main_rotater112_in[22], zll_main_rotater112_in[20], zll_main_rotater112_in[19], zll_main_rotater112_in[18], zll_main_rotater112_in[17], zll_main_rotater112_in[16], zll_main_rotater112_in[15], zll_main_rotater112_in[14], zll_main_rotater112_in[13], zll_main_rotater112_in[12], zll_main_rotater112_in[11], zll_main_rotater112_in[10], zll_main_rotater112_in[9], zll_main_rotater112_in[8], zll_main_rotater112_in[7], zll_main_rotater112_in[6], zll_main_rotater112_in[5], zll_main_rotater112_in[4], zll_main_rotater112_in[3], zll_main_rotater112_in[2], zll_main_rotater112_in[1], zll_main_rotater112_in[0]};
  assign zll_main_rotater1130_in = {zll_main_rotater1119_in[31], zll_main_rotater1119_in[30], zll_main_rotater1119_in[29], zll_main_rotater1119_in[28], zll_main_rotater1119_in[27], zll_main_rotater1119_in[26], zll_main_rotater1119_in[25], zll_main_rotater1119_in[24], zll_main_rotater1119_in[20], zll_main_rotater1119_in[23], zll_main_rotater1119_in[22], zll_main_rotater1119_in[21], zll_main_rotater1119_in[19], zll_main_rotater1119_in[18], zll_main_rotater1119_in[17], zll_main_rotater1119_in[16], zll_main_rotater1119_in[15], zll_main_rotater1119_in[14], zll_main_rotater1119_in[13], zll_main_rotater1119_in[12], zll_main_rotater1119_in[11], zll_main_rotater1119_in[10], zll_main_rotater1119_in[9], zll_main_rotater1119_in[8], zll_main_rotater1119_in[7], zll_main_rotater1119_in[6], zll_main_rotater1119_in[5], zll_main_rotater1119_in[4], zll_main_rotater1119_in[3], zll_main_rotater1119_in[2], zll_main_rotater1119_in[1], zll_main_rotater1119_in[0]};
  assign zll_main_rotater111_in = {zll_main_rotater1130_in[31], zll_main_rotater1130_in[30], zll_main_rotater1130_in[29], zll_main_rotater1130_in[28], zll_main_rotater1130_in[27], zll_main_rotater1130_in[19], zll_main_rotater1130_in[26], zll_main_rotater1130_in[25], zll_main_rotater1130_in[24], zll_main_rotater1130_in[23], zll_main_rotater1130_in[22], zll_main_rotater1130_in[21], zll_main_rotater1130_in[20], zll_main_rotater1130_in[18], zll_main_rotater1130_in[17], zll_main_rotater1130_in[16], zll_main_rotater1130_in[15], zll_main_rotater1130_in[14], zll_main_rotater1130_in[13], zll_main_rotater1130_in[12], zll_main_rotater1130_in[11], zll_main_rotater1130_in[10], zll_main_rotater1130_in[9], zll_main_rotater1130_in[8], zll_main_rotater1130_in[7], zll_main_rotater1130_in[6], zll_main_rotater1130_in[5], zll_main_rotater1130_in[4], zll_main_rotater1130_in[3], zll_main_rotater1130_in[2], zll_main_rotater1130_in[1], zll_main_rotater1130_in[0]};
  assign zll_main_rotater1111_in = {zll_main_rotater111_in[31], zll_main_rotater111_in[30], zll_main_rotater111_in[29], zll_main_rotater111_in[28], zll_main_rotater111_in[27], zll_main_rotater111_in[26], zll_main_rotater111_in[25], zll_main_rotater111_in[24], zll_main_rotater111_in[23], zll_main_rotater111_in[22], zll_main_rotater111_in[18], zll_main_rotater111_in[21], zll_main_rotater111_in[20], zll_main_rotater111_in[19], zll_main_rotater111_in[17], zll_main_rotater111_in[16], zll_main_rotater111_in[15], zll_main_rotater111_in[14], zll_main_rotater111_in[13], zll_main_rotater111_in[12], zll_main_rotater111_in[11], zll_main_rotater111_in[10], zll_main_rotater111_in[9], zll_main_rotater111_in[8], zll_main_rotater111_in[7], zll_main_rotater111_in[6], zll_main_rotater111_in[5], zll_main_rotater111_in[4], zll_main_rotater111_in[3], zll_main_rotater111_in[2], zll_main_rotater111_in[1], zll_main_rotater111_in[0]};
  assign zll_main_rotater119_in = {zll_main_rotater1111_in[31], zll_main_rotater1111_in[30], zll_main_rotater1111_in[17], zll_main_rotater1111_in[29], zll_main_rotater1111_in[28], zll_main_rotater1111_in[27], zll_main_rotater1111_in[26], zll_main_rotater1111_in[25], zll_main_rotater1111_in[24], zll_main_rotater1111_in[23], zll_main_rotater1111_in[22], zll_main_rotater1111_in[21], zll_main_rotater1111_in[20], zll_main_rotater1111_in[19], zll_main_rotater1111_in[18], zll_main_rotater1111_in[16], zll_main_rotater1111_in[15], zll_main_rotater1111_in[14], zll_main_rotater1111_in[13], zll_main_rotater1111_in[12], zll_main_rotater1111_in[11], zll_main_rotater1111_in[10], zll_main_rotater1111_in[9], zll_main_rotater1111_in[8], zll_main_rotater1111_in[7], zll_main_rotater1111_in[6], zll_main_rotater1111_in[5], zll_main_rotater1111_in[4], zll_main_rotater1111_in[3], zll_main_rotater1111_in[2], zll_main_rotater1111_in[1], zll_main_rotater1111_in[0]};
  assign zll_main_rotater1125_in = {zll_main_rotater119_in[16], zll_main_rotater119_in[31], zll_main_rotater119_in[30], zll_main_rotater119_in[29], zll_main_rotater119_in[28], zll_main_rotater119_in[27], zll_main_rotater119_in[26], zll_main_rotater119_in[25], zll_main_rotater119_in[24], zll_main_rotater119_in[23], zll_main_rotater119_in[22], zll_main_rotater119_in[21], zll_main_rotater119_in[20], zll_main_rotater119_in[19], zll_main_rotater119_in[18], zll_main_rotater119_in[17], zll_main_rotater119_in[15], zll_main_rotater119_in[14], zll_main_rotater119_in[13], zll_main_rotater119_in[12], zll_main_rotater119_in[11], zll_main_rotater119_in[10], zll_main_rotater119_in[9], zll_main_rotater119_in[8], zll_main_rotater119_in[7], zll_main_rotater119_in[6], zll_main_rotater119_in[5], zll_main_rotater119_in[4], zll_main_rotater119_in[3], zll_main_rotater119_in[2], zll_main_rotater119_in[1], zll_main_rotater119_in[0]};
  assign zll_main_rotater1127_in = {zll_main_rotater1125_in[31], zll_main_rotater1125_in[30], zll_main_rotater1125_in[29], zll_main_rotater1125_in[28], zll_main_rotater1125_in[27], zll_main_rotater1125_in[26], zll_main_rotater1125_in[25], zll_main_rotater1125_in[24], zll_main_rotater1125_in[23], zll_main_rotater1125_in[15], zll_main_rotater1125_in[22], zll_main_rotater1125_in[21], zll_main_rotater1125_in[20], zll_main_rotater1125_in[19], zll_main_rotater1125_in[18], zll_main_rotater1125_in[17], zll_main_rotater1125_in[16], zll_main_rotater1125_in[14], zll_main_rotater1125_in[13], zll_main_rotater1125_in[12], zll_main_rotater1125_in[11], zll_main_rotater1125_in[10], zll_main_rotater1125_in[9], zll_main_rotater1125_in[8], zll_main_rotater1125_in[7], zll_main_rotater1125_in[6], zll_main_rotater1125_in[5], zll_main_rotater1125_in[4], zll_main_rotater1125_in[3], zll_main_rotater1125_in[2], zll_main_rotater1125_in[1], zll_main_rotater1125_in[0]};
  assign zll_main_rotater1113_in = {zll_main_rotater1127_in[31], zll_main_rotater1127_in[30], zll_main_rotater1127_in[29], zll_main_rotater1127_in[28], zll_main_rotater1127_in[27], zll_main_rotater1127_in[26], zll_main_rotater1127_in[25], zll_main_rotater1127_in[24], zll_main_rotater1127_in[23], zll_main_rotater1127_in[22], zll_main_rotater1127_in[21], zll_main_rotater1127_in[20], zll_main_rotater1127_in[14], zll_main_rotater1127_in[19], zll_main_rotater1127_in[18], zll_main_rotater1127_in[17], zll_main_rotater1127_in[16], zll_main_rotater1127_in[15], zll_main_rotater1127_in[13], zll_main_rotater1127_in[12], zll_main_rotater1127_in[11], zll_main_rotater1127_in[10], zll_main_rotater1127_in[9], zll_main_rotater1127_in[8], zll_main_rotater1127_in[7], zll_main_rotater1127_in[6], zll_main_rotater1127_in[5], zll_main_rotater1127_in[4], zll_main_rotater1127_in[3], zll_main_rotater1127_in[2], zll_main_rotater1127_in[1], zll_main_rotater1127_in[0]};
  assign zll_main_rotater1128_in = {zll_main_rotater1113_in[31], zll_main_rotater1113_in[30], zll_main_rotater1113_in[29], zll_main_rotater1113_in[28], zll_main_rotater1113_in[27], zll_main_rotater1113_in[26], zll_main_rotater1113_in[13], zll_main_rotater1113_in[25], zll_main_rotater1113_in[24], zll_main_rotater1113_in[23], zll_main_rotater1113_in[22], zll_main_rotater1113_in[21], zll_main_rotater1113_in[20], zll_main_rotater1113_in[19], zll_main_rotater1113_in[18], zll_main_rotater1113_in[17], zll_main_rotater1113_in[16], zll_main_rotater1113_in[15], zll_main_rotater1113_in[14], zll_main_rotater1113_in[12], zll_main_rotater1113_in[11], zll_main_rotater1113_in[10], zll_main_rotater1113_in[9], zll_main_rotater1113_in[8], zll_main_rotater1113_in[7], zll_main_rotater1113_in[6], zll_main_rotater1113_in[5], zll_main_rotater1113_in[4], zll_main_rotater1113_in[3], zll_main_rotater1113_in[2], zll_main_rotater1113_in[1], zll_main_rotater1113_in[0]};
  assign zll_main_rotater11_in = {zll_main_rotater1128_in[31], zll_main_rotater1128_in[30], zll_main_rotater1128_in[29], zll_main_rotater1128_in[28], zll_main_rotater1128_in[27], zll_main_rotater1128_in[26], zll_main_rotater1128_in[25], zll_main_rotater1128_in[24], zll_main_rotater1128_in[23], zll_main_rotater1128_in[22], zll_main_rotater1128_in[21], zll_main_rotater1128_in[20], zll_main_rotater1128_in[12], zll_main_rotater1128_in[19], zll_main_rotater1128_in[18], zll_main_rotater1128_in[17], zll_main_rotater1128_in[16], zll_main_rotater1128_in[15], zll_main_rotater1128_in[14], zll_main_rotater1128_in[13], zll_main_rotater1128_in[11], zll_main_rotater1128_in[10], zll_main_rotater1128_in[9], zll_main_rotater1128_in[8], zll_main_rotater1128_in[7], zll_main_rotater1128_in[6], zll_main_rotater1128_in[5], zll_main_rotater1128_in[4], zll_main_rotater1128_in[3], zll_main_rotater1128_in[2], zll_main_rotater1128_in[1], zll_main_rotater1128_in[0]};
  assign zll_main_rotater1118_in = {zll_main_rotater11_in[31], zll_main_rotater11_in[30], zll_main_rotater11_in[29], zll_main_rotater11_in[28], zll_main_rotater11_in[27], zll_main_rotater11_in[26], zll_main_rotater11_in[25], zll_main_rotater11_in[24], zll_main_rotater11_in[23], zll_main_rotater11_in[22], zll_main_rotater11_in[21], zll_main_rotater11_in[20], zll_main_rotater11_in[19], zll_main_rotater11_in[18], zll_main_rotater11_in[17], zll_main_rotater11_in[16], zll_main_rotater11_in[11], zll_main_rotater11_in[15], zll_main_rotater11_in[14], zll_main_rotater11_in[13], zll_main_rotater11_in[12], zll_main_rotater11_in[10], zll_main_rotater11_in[9], zll_main_rotater11_in[8], zll_main_rotater11_in[7], zll_main_rotater11_in[6], zll_main_rotater11_in[5], zll_main_rotater11_in[4], zll_main_rotater11_in[3], zll_main_rotater11_in[2], zll_main_rotater11_in[1], zll_main_rotater11_in[0]};
  assign zll_main_rotater1114_in = {zll_main_rotater1118_in[31], zll_main_rotater1118_in[30], zll_main_rotater1118_in[29], zll_main_rotater1118_in[28], zll_main_rotater1118_in[27], zll_main_rotater1118_in[26], zll_main_rotater1118_in[25], zll_main_rotater1118_in[24], zll_main_rotater1118_in[23], zll_main_rotater1118_in[22], zll_main_rotater1118_in[21], zll_main_rotater1118_in[20], zll_main_rotater1118_in[19], zll_main_rotater1118_in[18], zll_main_rotater1118_in[17], zll_main_rotater1118_in[16], zll_main_rotater1118_in[15], zll_main_rotater1118_in[14], zll_main_rotater1118_in[13], zll_main_rotater1118_in[10], zll_main_rotater1118_in[12], zll_main_rotater1118_in[11], zll_main_rotater1118_in[9], zll_main_rotater1118_in[8], zll_main_rotater1118_in[7], zll_main_rotater1118_in[6], zll_main_rotater1118_in[5], zll_main_rotater1118_in[4], zll_main_rotater1118_in[3], zll_main_rotater1118_in[2], zll_main_rotater1118_in[1], zll_main_rotater1118_in[0]};
  assign zll_main_rotater117_in = {zll_main_rotater1114_in[31], zll_main_rotater1114_in[30], zll_main_rotater1114_in[29], zll_main_rotater1114_in[28], zll_main_rotater1114_in[27], zll_main_rotater1114_in[26], zll_main_rotater1114_in[25], zll_main_rotater1114_in[24], zll_main_rotater1114_in[23], zll_main_rotater1114_in[22], zll_main_rotater1114_in[21], zll_main_rotater1114_in[20], zll_main_rotater1114_in[19], zll_main_rotater1114_in[18], zll_main_rotater1114_in[17], zll_main_rotater1114_in[16], zll_main_rotater1114_in[15], zll_main_rotater1114_in[14], zll_main_rotater1114_in[13], zll_main_rotater1114_in[12], zll_main_rotater1114_in[11], zll_main_rotater1114_in[9], zll_main_rotater1114_in[10], zll_main_rotater1114_in[8], zll_main_rotater1114_in[7], zll_main_rotater1114_in[6], zll_main_rotater1114_in[5], zll_main_rotater1114_in[4], zll_main_rotater1114_in[3], zll_main_rotater1114_in[2], zll_main_rotater1114_in[1], zll_main_rotater1114_in[0]};
  assign zll_main_rotater1115_in = {zll_main_rotater117_in[31], zll_main_rotater117_in[30], zll_main_rotater117_in[29], zll_main_rotater117_in[28], zll_main_rotater117_in[27], zll_main_rotater117_in[26], zll_main_rotater117_in[25], zll_main_rotater117_in[24], zll_main_rotater117_in[23], zll_main_rotater117_in[22], zll_main_rotater117_in[21], zll_main_rotater117_in[20], zll_main_rotater117_in[19], zll_main_rotater117_in[8], zll_main_rotater117_in[18], zll_main_rotater117_in[17], zll_main_rotater117_in[16], zll_main_rotater117_in[15], zll_main_rotater117_in[14], zll_main_rotater117_in[13], zll_main_rotater117_in[12], zll_main_rotater117_in[11], zll_main_rotater117_in[10], zll_main_rotater117_in[9], zll_main_rotater117_in[7], zll_main_rotater117_in[6], zll_main_rotater117_in[5], zll_main_rotater117_in[4], zll_main_rotater117_in[3], zll_main_rotater117_in[2], zll_main_rotater117_in[1], zll_main_rotater117_in[0]};
  assign zll_main_rotater1116_in = {zll_main_rotater1115_in[31], zll_main_rotater1115_in[30], zll_main_rotater1115_in[29], zll_main_rotater1115_in[28], zll_main_rotater1115_in[27], zll_main_rotater1115_in[26], zll_main_rotater1115_in[25], zll_main_rotater1115_in[24], zll_main_rotater1115_in[7], zll_main_rotater1115_in[23], zll_main_rotater1115_in[22], zll_main_rotater1115_in[21], zll_main_rotater1115_in[20], zll_main_rotater1115_in[19], zll_main_rotater1115_in[18], zll_main_rotater1115_in[17], zll_main_rotater1115_in[16], zll_main_rotater1115_in[15], zll_main_rotater1115_in[14], zll_main_rotater1115_in[13], zll_main_rotater1115_in[12], zll_main_rotater1115_in[11], zll_main_rotater1115_in[10], zll_main_rotater1115_in[9], zll_main_rotater1115_in[8], zll_main_rotater1115_in[6], zll_main_rotater1115_in[5], zll_main_rotater1115_in[4], zll_main_rotater1115_in[3], zll_main_rotater1115_in[2], zll_main_rotater1115_in[1], zll_main_rotater1115_in[0]};
  assign zll_main_rotater113_in = {zll_main_rotater1116_in[6], zll_main_rotater1116_in[31], zll_main_rotater1116_in[30], zll_main_rotater1116_in[29], zll_main_rotater1116_in[28], zll_main_rotater1116_in[27], zll_main_rotater1116_in[26], zll_main_rotater1116_in[25], zll_main_rotater1116_in[24], zll_main_rotater1116_in[23], zll_main_rotater1116_in[22], zll_main_rotater1116_in[21], zll_main_rotater1116_in[20], zll_main_rotater1116_in[19], zll_main_rotater1116_in[18], zll_main_rotater1116_in[17], zll_main_rotater1116_in[16], zll_main_rotater1116_in[15], zll_main_rotater1116_in[14], zll_main_rotater1116_in[13], zll_main_rotater1116_in[12], zll_main_rotater1116_in[11], zll_main_rotater1116_in[10], zll_main_rotater1116_in[9], zll_main_rotater1116_in[8], zll_main_rotater1116_in[7], zll_main_rotater1116_in[5], zll_main_rotater1116_in[4], zll_main_rotater1116_in[3], zll_main_rotater1116_in[2], zll_main_rotater1116_in[1], zll_main_rotater1116_in[0]};
  assign zll_main_rotater115_in = {zll_main_rotater113_in[31], zll_main_rotater113_in[30], zll_main_rotater113_in[29], zll_main_rotater113_in[28], zll_main_rotater113_in[27], zll_main_rotater113_in[26], zll_main_rotater113_in[25], zll_main_rotater113_in[24], zll_main_rotater113_in[23], zll_main_rotater113_in[22], zll_main_rotater113_in[21], zll_main_rotater113_in[20], zll_main_rotater113_in[19], zll_main_rotater113_in[18], zll_main_rotater113_in[17], zll_main_rotater113_in[16], zll_main_rotater113_in[15], zll_main_rotater113_in[14], zll_main_rotater113_in[13], zll_main_rotater113_in[5], zll_main_rotater113_in[12], zll_main_rotater113_in[11], zll_main_rotater113_in[10], zll_main_rotater113_in[9], zll_main_rotater113_in[8], zll_main_rotater113_in[7], zll_main_rotater113_in[6], zll_main_rotater113_in[4], zll_main_rotater113_in[3], zll_main_rotater113_in[2], zll_main_rotater113_in[1], zll_main_rotater113_in[0]};
  assign zll_main_rotater1112_in = {zll_main_rotater115_in[31], zll_main_rotater115_in[30], zll_main_rotater115_in[29], zll_main_rotater115_in[28], zll_main_rotater115_in[27], zll_main_rotater115_in[26], zll_main_rotater115_in[25], zll_main_rotater115_in[24], zll_main_rotater115_in[23], zll_main_rotater115_in[22], zll_main_rotater115_in[21], zll_main_rotater115_in[20], zll_main_rotater115_in[19], zll_main_rotater115_in[18], zll_main_rotater115_in[17], zll_main_rotater115_in[16], zll_main_rotater115_in[15], zll_main_rotater115_in[14], zll_main_rotater115_in[13], zll_main_rotater115_in[4], zll_main_rotater115_in[12], zll_main_rotater115_in[11], zll_main_rotater115_in[10], zll_main_rotater115_in[9], zll_main_rotater115_in[8], zll_main_rotater115_in[7], zll_main_rotater115_in[6], zll_main_rotater115_in[5], zll_main_rotater115_in[3], zll_main_rotater115_in[2], zll_main_rotater115_in[1], zll_main_rotater115_in[0]};
  assign zll_main_rotater1120_in = {zll_main_rotater1112_in[31], zll_main_rotater1112_in[30], zll_main_rotater1112_in[29], zll_main_rotater1112_in[28], zll_main_rotater1112_in[27], zll_main_rotater1112_in[26], zll_main_rotater1112_in[25], zll_main_rotater1112_in[24], zll_main_rotater1112_in[23], zll_main_rotater1112_in[22], zll_main_rotater1112_in[21], zll_main_rotater1112_in[3], zll_main_rotater1112_in[20], zll_main_rotater1112_in[19], zll_main_rotater1112_in[18], zll_main_rotater1112_in[17], zll_main_rotater1112_in[16], zll_main_rotater1112_in[15], zll_main_rotater1112_in[14], zll_main_rotater1112_in[13], zll_main_rotater1112_in[12], zll_main_rotater1112_in[11], zll_main_rotater1112_in[10], zll_main_rotater1112_in[9], zll_main_rotater1112_in[8], zll_main_rotater1112_in[7], zll_main_rotater1112_in[6], zll_main_rotater1112_in[5], zll_main_rotater1112_in[4], zll_main_rotater1112_in[2], zll_main_rotater1112_in[1], zll_main_rotater1112_in[0]};
  assign zll_main_rotater1131_in = {zll_main_rotater1120_in[2], zll_main_rotater1120_in[31], zll_main_rotater1120_in[30], zll_main_rotater1120_in[29], zll_main_rotater1120_in[28], zll_main_rotater1120_in[27], zll_main_rotater1120_in[26], zll_main_rotater1120_in[25], zll_main_rotater1120_in[24], zll_main_rotater1120_in[23], zll_main_rotater1120_in[22], zll_main_rotater1120_in[21], zll_main_rotater1120_in[20], zll_main_rotater1120_in[19], zll_main_rotater1120_in[18], zll_main_rotater1120_in[17], zll_main_rotater1120_in[16], zll_main_rotater1120_in[15], zll_main_rotater1120_in[14], zll_main_rotater1120_in[13], zll_main_rotater1120_in[12], zll_main_rotater1120_in[11], zll_main_rotater1120_in[10], zll_main_rotater1120_in[9], zll_main_rotater1120_in[8], zll_main_rotater1120_in[7], zll_main_rotater1120_in[6], zll_main_rotater1120_in[5], zll_main_rotater1120_in[4], zll_main_rotater1120_in[3], zll_main_rotater1120_in[1], zll_main_rotater1120_in[0]};
  assign xorw32_in = {{zll_main_rotater626_in[28], zll_main_rotater626_in[22], zll_main_rotater626_in[4], zll_main_rotater626_in[25], zll_main_rotater626_in[16], zll_main_rotater626_in[0], zll_main_rotater626_in[3], zll_main_rotater626_in[17], zll_main_rotater626_in[18], zll_main_rotater626_in[2], zll_main_rotater626_in[21], zll_main_rotater626_in[27], zll_main_rotater626_in[7], zll_main_rotater626_in[14], zll_main_rotater626_in[8], zll_main_rotater626_in[10], zll_main_rotater626_in[15], zll_main_rotater626_in[12], zll_main_rotater626_in[1], zll_main_rotater626_in[23], zll_main_rotater626_in[20], zll_main_rotater626_in[9], zll_main_rotater626_in[24], zll_main_rotater626_in[11], zll_main_rotater626_in[13], zll_main_rotater626_in[5], zll_main_rotater626_in[19], zll_main_rotater626_in[31], zll_main_rotater626_in[30], zll_main_rotater626_in[6], zll_main_rotater626_in[26], zll_main_rotater626_in[29]}, {zll_main_rotater1131_in[5], zll_main_rotater1131_in[3], zll_main_rotater1131_in[14], zll_main_rotater1131_in[21], zll_main_rotater1131_in[30], zll_main_rotater1131_in[9], zll_main_rotater1131_in[10], zll_main_rotater1131_in[19], zll_main_rotater1131_in[31], zll_main_rotater1131_in[1], zll_main_rotater1131_in[0], zll_main_rotater1131_in[24], zll_main_rotater1131_in[16], zll_main_rotater1131_in[22], zll_main_rotater1131_in[25], zll_main_rotater1131_in[18], zll_main_rotater1131_in[13], zll_main_rotater1131_in[4], zll_main_rotater1131_in[27], zll_main_rotater1131_in[28], zll_main_rotater1131_in[2], zll_main_rotater1131_in[6], zll_main_rotater1131_in[11], zll_main_rotater1131_in[20], zll_main_rotater1131_in[7], zll_main_rotater1131_in[26], zll_main_rotater1131_in[29], zll_main_rotater1131_in[17], zll_main_rotater1131_in[12], zll_main_rotater1131_in[23], zll_main_rotater1131_in[15], zll_main_rotater1131_in[8]}};
  xorW32  inst (xorw32_in[63:32], xorw32_in[31:0], extres[31:0]);
  assign main_rotater25_in = arg0;
  assign zll_main_rotater2521_in = main_rotater25_in[31:0];
  assign zll_main_rotater2515_in = {zll_main_rotater2521_in[31], zll_main_rotater2521_in[30], zll_main_rotater2521_in[28], zll_main_rotater2521_in[29], zll_main_rotater2521_in[27], zll_main_rotater2521_in[26], zll_main_rotater2521_in[25], zll_main_rotater2521_in[24], zll_main_rotater2521_in[23], zll_main_rotater2521_in[22], zll_main_rotater2521_in[21], zll_main_rotater2521_in[20], zll_main_rotater2521_in[19], zll_main_rotater2521_in[18], zll_main_rotater2521_in[17], zll_main_rotater2521_in[16], zll_main_rotater2521_in[15], zll_main_rotater2521_in[14], zll_main_rotater2521_in[13], zll_main_rotater2521_in[12], zll_main_rotater2521_in[11], zll_main_rotater2521_in[10], zll_main_rotater2521_in[9], zll_main_rotater2521_in[8], zll_main_rotater2521_in[7], zll_main_rotater2521_in[6], zll_main_rotater2521_in[5], zll_main_rotater2521_in[4], zll_main_rotater2521_in[3], zll_main_rotater2521_in[2], zll_main_rotater2521_in[1], zll_main_rotater2521_in[0]};
  assign zll_main_rotater2518_in = {zll_main_rotater2515_in[31], zll_main_rotater2515_in[30], zll_main_rotater2515_in[29], zll_main_rotater2515_in[27], zll_main_rotater2515_in[28], zll_main_rotater2515_in[26], zll_main_rotater2515_in[25], zll_main_rotater2515_in[24], zll_main_rotater2515_in[23], zll_main_rotater2515_in[22], zll_main_rotater2515_in[21], zll_main_rotater2515_in[20], zll_main_rotater2515_in[19], zll_main_rotater2515_in[18], zll_main_rotater2515_in[17], zll_main_rotater2515_in[16], zll_main_rotater2515_in[15], zll_main_rotater2515_in[14], zll_main_rotater2515_in[13], zll_main_rotater2515_in[12], zll_main_rotater2515_in[11], zll_main_rotater2515_in[10], zll_main_rotater2515_in[9], zll_main_rotater2515_in[8], zll_main_rotater2515_in[7], zll_main_rotater2515_in[6], zll_main_rotater2515_in[5], zll_main_rotater2515_in[4], zll_main_rotater2515_in[3], zll_main_rotater2515_in[2], zll_main_rotater2515_in[1], zll_main_rotater2515_in[0]};
  assign zll_main_rotater2516_in = {zll_main_rotater2518_in[31], zll_main_rotater2518_in[26], zll_main_rotater2518_in[30], zll_main_rotater2518_in[29], zll_main_rotater2518_in[28], zll_main_rotater2518_in[27], zll_main_rotater2518_in[25], zll_main_rotater2518_in[24], zll_main_rotater2518_in[23], zll_main_rotater2518_in[22], zll_main_rotater2518_in[21], zll_main_rotater2518_in[20], zll_main_rotater2518_in[19], zll_main_rotater2518_in[18], zll_main_rotater2518_in[17], zll_main_rotater2518_in[16], zll_main_rotater2518_in[15], zll_main_rotater2518_in[14], zll_main_rotater2518_in[13], zll_main_rotater2518_in[12], zll_main_rotater2518_in[11], zll_main_rotater2518_in[10], zll_main_rotater2518_in[9], zll_main_rotater2518_in[8], zll_main_rotater2518_in[7], zll_main_rotater2518_in[6], zll_main_rotater2518_in[5], zll_main_rotater2518_in[4], zll_main_rotater2518_in[3], zll_main_rotater2518_in[2], zll_main_rotater2518_in[1], zll_main_rotater2518_in[0]};
  assign zll_main_rotater251_in = {zll_main_rotater2516_in[31], zll_main_rotater2516_in[30], zll_main_rotater2516_in[29], zll_main_rotater2516_in[28], zll_main_rotater2516_in[27], zll_main_rotater2516_in[25], zll_main_rotater2516_in[26], zll_main_rotater2516_in[24], zll_main_rotater2516_in[23], zll_main_rotater2516_in[22], zll_main_rotater2516_in[21], zll_main_rotater2516_in[20], zll_main_rotater2516_in[19], zll_main_rotater2516_in[18], zll_main_rotater2516_in[17], zll_main_rotater2516_in[16], zll_main_rotater2516_in[15], zll_main_rotater2516_in[14], zll_main_rotater2516_in[13], zll_main_rotater2516_in[12], zll_main_rotater2516_in[11], zll_main_rotater2516_in[10], zll_main_rotater2516_in[9], zll_main_rotater2516_in[8], zll_main_rotater2516_in[7], zll_main_rotater2516_in[6], zll_main_rotater2516_in[5], zll_main_rotater2516_in[4], zll_main_rotater2516_in[3], zll_main_rotater2516_in[2], zll_main_rotater2516_in[1], zll_main_rotater2516_in[0]};
  assign zll_main_rotater2526_in = {zll_main_rotater251_in[31], zll_main_rotater251_in[30], zll_main_rotater251_in[29], zll_main_rotater251_in[28], zll_main_rotater251_in[24], zll_main_rotater251_in[27], zll_main_rotater251_in[26], zll_main_rotater251_in[25], zll_main_rotater251_in[23], zll_main_rotater251_in[22], zll_main_rotater251_in[21], zll_main_rotater251_in[20], zll_main_rotater251_in[19], zll_main_rotater251_in[18], zll_main_rotater251_in[17], zll_main_rotater251_in[16], zll_main_rotater251_in[15], zll_main_rotater251_in[14], zll_main_rotater251_in[13], zll_main_rotater251_in[12], zll_main_rotater251_in[11], zll_main_rotater251_in[10], zll_main_rotater251_in[9], zll_main_rotater251_in[8], zll_main_rotater251_in[7], zll_main_rotater251_in[6], zll_main_rotater251_in[5], zll_main_rotater251_in[4], zll_main_rotater251_in[3], zll_main_rotater251_in[2], zll_main_rotater251_in[1], zll_main_rotater251_in[0]};
  assign zll_main_rotater255_in = {zll_main_rotater2526_in[31], zll_main_rotater2526_in[30], zll_main_rotater2526_in[29], zll_main_rotater2526_in[28], zll_main_rotater2526_in[23], zll_main_rotater2526_in[27], zll_main_rotater2526_in[26], zll_main_rotater2526_in[25], zll_main_rotater2526_in[24], zll_main_rotater2526_in[22], zll_main_rotater2526_in[21], zll_main_rotater2526_in[20], zll_main_rotater2526_in[19], zll_main_rotater2526_in[18], zll_main_rotater2526_in[17], zll_main_rotater2526_in[16], zll_main_rotater2526_in[15], zll_main_rotater2526_in[14], zll_main_rotater2526_in[13], zll_main_rotater2526_in[12], zll_main_rotater2526_in[11], zll_main_rotater2526_in[10], zll_main_rotater2526_in[9], zll_main_rotater2526_in[8], zll_main_rotater2526_in[7], zll_main_rotater2526_in[6], zll_main_rotater2526_in[5], zll_main_rotater2526_in[4], zll_main_rotater2526_in[3], zll_main_rotater2526_in[2], zll_main_rotater2526_in[1], zll_main_rotater2526_in[0]};
  assign zll_main_rotater2528_in = {zll_main_rotater255_in[31], zll_main_rotater255_in[30], zll_main_rotater255_in[29], zll_main_rotater255_in[28], zll_main_rotater255_in[27], zll_main_rotater255_in[26], zll_main_rotater255_in[25], zll_main_rotater255_in[24], zll_main_rotater255_in[22], zll_main_rotater255_in[23], zll_main_rotater255_in[21], zll_main_rotater255_in[20], zll_main_rotater255_in[19], zll_main_rotater255_in[18], zll_main_rotater255_in[17], zll_main_rotater255_in[16], zll_main_rotater255_in[15], zll_main_rotater255_in[14], zll_main_rotater255_in[13], zll_main_rotater255_in[12], zll_main_rotater255_in[11], zll_main_rotater255_in[10], zll_main_rotater255_in[9], zll_main_rotater255_in[8], zll_main_rotater255_in[7], zll_main_rotater255_in[6], zll_main_rotater255_in[5], zll_main_rotater255_in[4], zll_main_rotater255_in[3], zll_main_rotater255_in[2], zll_main_rotater255_in[1], zll_main_rotater255_in[0]};
  assign zll_main_rotater2511_in = {zll_main_rotater2528_in[31], zll_main_rotater2528_in[21], zll_main_rotater2528_in[30], zll_main_rotater2528_in[29], zll_main_rotater2528_in[28], zll_main_rotater2528_in[27], zll_main_rotater2528_in[26], zll_main_rotater2528_in[25], zll_main_rotater2528_in[24], zll_main_rotater2528_in[23], zll_main_rotater2528_in[22], zll_main_rotater2528_in[20], zll_main_rotater2528_in[19], zll_main_rotater2528_in[18], zll_main_rotater2528_in[17], zll_main_rotater2528_in[16], zll_main_rotater2528_in[15], zll_main_rotater2528_in[14], zll_main_rotater2528_in[13], zll_main_rotater2528_in[12], zll_main_rotater2528_in[11], zll_main_rotater2528_in[10], zll_main_rotater2528_in[9], zll_main_rotater2528_in[8], zll_main_rotater2528_in[7], zll_main_rotater2528_in[6], zll_main_rotater2528_in[5], zll_main_rotater2528_in[4], zll_main_rotater2528_in[3], zll_main_rotater2528_in[2], zll_main_rotater2528_in[1], zll_main_rotater2528_in[0]};
  assign zll_main_rotater259_in = {zll_main_rotater2511_in[31], zll_main_rotater2511_in[19], zll_main_rotater2511_in[30], zll_main_rotater2511_in[29], zll_main_rotater2511_in[28], zll_main_rotater2511_in[27], zll_main_rotater2511_in[26], zll_main_rotater2511_in[25], zll_main_rotater2511_in[24], zll_main_rotater2511_in[23], zll_main_rotater2511_in[22], zll_main_rotater2511_in[21], zll_main_rotater2511_in[20], zll_main_rotater2511_in[18], zll_main_rotater2511_in[17], zll_main_rotater2511_in[16], zll_main_rotater2511_in[15], zll_main_rotater2511_in[14], zll_main_rotater2511_in[13], zll_main_rotater2511_in[12], zll_main_rotater2511_in[11], zll_main_rotater2511_in[10], zll_main_rotater2511_in[9], zll_main_rotater2511_in[8], zll_main_rotater2511_in[7], zll_main_rotater2511_in[6], zll_main_rotater2511_in[5], zll_main_rotater2511_in[4], zll_main_rotater2511_in[3], zll_main_rotater2511_in[2], zll_main_rotater2511_in[1], zll_main_rotater2511_in[0]};
  assign zll_main_rotater2510_in = {zll_main_rotater259_in[31], zll_main_rotater259_in[30], zll_main_rotater259_in[29], zll_main_rotater259_in[28], zll_main_rotater259_in[27], zll_main_rotater259_in[26], zll_main_rotater259_in[25], zll_main_rotater259_in[24], zll_main_rotater259_in[18], zll_main_rotater259_in[23], zll_main_rotater259_in[22], zll_main_rotater259_in[21], zll_main_rotater259_in[20], zll_main_rotater259_in[19], zll_main_rotater259_in[17], zll_main_rotater259_in[16], zll_main_rotater259_in[15], zll_main_rotater259_in[14], zll_main_rotater259_in[13], zll_main_rotater259_in[12], zll_main_rotater259_in[11], zll_main_rotater259_in[10], zll_main_rotater259_in[9], zll_main_rotater259_in[8], zll_main_rotater259_in[7], zll_main_rotater259_in[6], zll_main_rotater259_in[5], zll_main_rotater259_in[4], zll_main_rotater259_in[3], zll_main_rotater259_in[2], zll_main_rotater259_in[1], zll_main_rotater259_in[0]};
  assign zll_main_rotater2527_in = {zll_main_rotater2510_in[31], zll_main_rotater2510_in[30], zll_main_rotater2510_in[29], zll_main_rotater2510_in[28], zll_main_rotater2510_in[27], zll_main_rotater2510_in[26], zll_main_rotater2510_in[25], zll_main_rotater2510_in[24], zll_main_rotater2510_in[23], zll_main_rotater2510_in[22], zll_main_rotater2510_in[21], zll_main_rotater2510_in[17], zll_main_rotater2510_in[20], zll_main_rotater2510_in[19], zll_main_rotater2510_in[18], zll_main_rotater2510_in[16], zll_main_rotater2510_in[15], zll_main_rotater2510_in[14], zll_main_rotater2510_in[13], zll_main_rotater2510_in[12], zll_main_rotater2510_in[11], zll_main_rotater2510_in[10], zll_main_rotater2510_in[9], zll_main_rotater2510_in[8], zll_main_rotater2510_in[7], zll_main_rotater2510_in[6], zll_main_rotater2510_in[5], zll_main_rotater2510_in[4], zll_main_rotater2510_in[3], zll_main_rotater2510_in[2], zll_main_rotater2510_in[1], zll_main_rotater2510_in[0]};
  assign zll_main_rotater2525_in = {zll_main_rotater2527_in[31], zll_main_rotater2527_in[30], zll_main_rotater2527_in[29], zll_main_rotater2527_in[15], zll_main_rotater2527_in[28], zll_main_rotater2527_in[27], zll_main_rotater2527_in[26], zll_main_rotater2527_in[25], zll_main_rotater2527_in[24], zll_main_rotater2527_in[23], zll_main_rotater2527_in[22], zll_main_rotater2527_in[21], zll_main_rotater2527_in[20], zll_main_rotater2527_in[19], zll_main_rotater2527_in[18], zll_main_rotater2527_in[17], zll_main_rotater2527_in[16], zll_main_rotater2527_in[14], zll_main_rotater2527_in[13], zll_main_rotater2527_in[12], zll_main_rotater2527_in[11], zll_main_rotater2527_in[10], zll_main_rotater2527_in[9], zll_main_rotater2527_in[8], zll_main_rotater2527_in[7], zll_main_rotater2527_in[6], zll_main_rotater2527_in[5], zll_main_rotater2527_in[4], zll_main_rotater2527_in[3], zll_main_rotater2527_in[2], zll_main_rotater2527_in[1], zll_main_rotater2527_in[0]};
  assign zll_main_rotater2520_in = {zll_main_rotater2525_in[31], zll_main_rotater2525_in[30], zll_main_rotater2525_in[29], zll_main_rotater2525_in[28], zll_main_rotater2525_in[27], zll_main_rotater2525_in[26], zll_main_rotater2525_in[25], zll_main_rotater2525_in[14], zll_main_rotater2525_in[24], zll_main_rotater2525_in[23], zll_main_rotater2525_in[22], zll_main_rotater2525_in[21], zll_main_rotater2525_in[20], zll_main_rotater2525_in[19], zll_main_rotater2525_in[18], zll_main_rotater2525_in[17], zll_main_rotater2525_in[16], zll_main_rotater2525_in[15], zll_main_rotater2525_in[13], zll_main_rotater2525_in[12], zll_main_rotater2525_in[11], zll_main_rotater2525_in[10], zll_main_rotater2525_in[9], zll_main_rotater2525_in[8], zll_main_rotater2525_in[7], zll_main_rotater2525_in[6], zll_main_rotater2525_in[5], zll_main_rotater2525_in[4], zll_main_rotater2525_in[3], zll_main_rotater2525_in[2], zll_main_rotater2525_in[1], zll_main_rotater2525_in[0]};
  assign zll_main_rotater2512_in = {zll_main_rotater2520_in[31], zll_main_rotater2520_in[30], zll_main_rotater2520_in[29], zll_main_rotater2520_in[28], zll_main_rotater2520_in[27], zll_main_rotater2520_in[26], zll_main_rotater2520_in[25], zll_main_rotater2520_in[24], zll_main_rotater2520_in[23], zll_main_rotater2520_in[22], zll_main_rotater2520_in[21], zll_main_rotater2520_in[20], zll_main_rotater2520_in[19], zll_main_rotater2520_in[18], zll_main_rotater2520_in[17], zll_main_rotater2520_in[16], zll_main_rotater2520_in[13], zll_main_rotater2520_in[15], zll_main_rotater2520_in[14], zll_main_rotater2520_in[12], zll_main_rotater2520_in[11], zll_main_rotater2520_in[10], zll_main_rotater2520_in[9], zll_main_rotater2520_in[8], zll_main_rotater2520_in[7], zll_main_rotater2520_in[6], zll_main_rotater2520_in[5], zll_main_rotater2520_in[4], zll_main_rotater2520_in[3], zll_main_rotater2520_in[2], zll_main_rotater2520_in[1], zll_main_rotater2520_in[0]};
  assign zll_main_rotater258_in = {zll_main_rotater2512_in[12], zll_main_rotater2512_in[31], zll_main_rotater2512_in[30], zll_main_rotater2512_in[29], zll_main_rotater2512_in[28], zll_main_rotater2512_in[27], zll_main_rotater2512_in[26], zll_main_rotater2512_in[25], zll_main_rotater2512_in[24], zll_main_rotater2512_in[23], zll_main_rotater2512_in[22], zll_main_rotater2512_in[21], zll_main_rotater2512_in[20], zll_main_rotater2512_in[19], zll_main_rotater2512_in[18], zll_main_rotater2512_in[17], zll_main_rotater2512_in[16], zll_main_rotater2512_in[15], zll_main_rotater2512_in[14], zll_main_rotater2512_in[13], zll_main_rotater2512_in[11], zll_main_rotater2512_in[10], zll_main_rotater2512_in[9], zll_main_rotater2512_in[8], zll_main_rotater2512_in[7], zll_main_rotater2512_in[6], zll_main_rotater2512_in[5], zll_main_rotater2512_in[4], zll_main_rotater2512_in[3], zll_main_rotater2512_in[2], zll_main_rotater2512_in[1], zll_main_rotater2512_in[0]};
  assign zll_main_rotater254_in = {zll_main_rotater258_in[31], zll_main_rotater258_in[30], zll_main_rotater258_in[29], zll_main_rotater258_in[28], zll_main_rotater258_in[27], zll_main_rotater258_in[26], zll_main_rotater258_in[25], zll_main_rotater258_in[24], zll_main_rotater258_in[23], zll_main_rotater258_in[22], zll_main_rotater258_in[21], zll_main_rotater258_in[20], zll_main_rotater258_in[19], zll_main_rotater258_in[18], zll_main_rotater258_in[17], zll_main_rotater258_in[16], zll_main_rotater258_in[15], zll_main_rotater258_in[14], zll_main_rotater258_in[13], zll_main_rotater258_in[11], zll_main_rotater258_in[12], zll_main_rotater258_in[10], zll_main_rotater258_in[9], zll_main_rotater258_in[8], zll_main_rotater258_in[7], zll_main_rotater258_in[6], zll_main_rotater258_in[5], zll_main_rotater258_in[4], zll_main_rotater258_in[3], zll_main_rotater258_in[2], zll_main_rotater258_in[1], zll_main_rotater258_in[0]};
  assign zll_main_rotater256_in = {zll_main_rotater254_in[31], zll_main_rotater254_in[30], zll_main_rotater254_in[29], zll_main_rotater254_in[28], zll_main_rotater254_in[27], zll_main_rotater254_in[26], zll_main_rotater254_in[25], zll_main_rotater254_in[24], zll_main_rotater254_in[23], zll_main_rotater254_in[22], zll_main_rotater254_in[21], zll_main_rotater254_in[20], zll_main_rotater254_in[19], zll_main_rotater254_in[18], zll_main_rotater254_in[17], zll_main_rotater254_in[16], zll_main_rotater254_in[15], zll_main_rotater254_in[14], zll_main_rotater254_in[13], zll_main_rotater254_in[10], zll_main_rotater254_in[12], zll_main_rotater254_in[11], zll_main_rotater254_in[9], zll_main_rotater254_in[8], zll_main_rotater254_in[7], zll_main_rotater254_in[6], zll_main_rotater254_in[5], zll_main_rotater254_in[4], zll_main_rotater254_in[3], zll_main_rotater254_in[2], zll_main_rotater254_in[1], zll_main_rotater254_in[0]};
  assign zll_main_rotater253_in = {zll_main_rotater256_in[31], zll_main_rotater256_in[30], zll_main_rotater256_in[29], zll_main_rotater256_in[28], zll_main_rotater256_in[27], zll_main_rotater256_in[26], zll_main_rotater256_in[25], zll_main_rotater256_in[24], zll_main_rotater256_in[23], zll_main_rotater256_in[22], zll_main_rotater256_in[9], zll_main_rotater256_in[21], zll_main_rotater256_in[20], zll_main_rotater256_in[19], zll_main_rotater256_in[18], zll_main_rotater256_in[17], zll_main_rotater256_in[16], zll_main_rotater256_in[15], zll_main_rotater256_in[14], zll_main_rotater256_in[13], zll_main_rotater256_in[12], zll_main_rotater256_in[11], zll_main_rotater256_in[10], zll_main_rotater256_in[8], zll_main_rotater256_in[7], zll_main_rotater256_in[6], zll_main_rotater256_in[5], zll_main_rotater256_in[4], zll_main_rotater256_in[3], zll_main_rotater256_in[2], zll_main_rotater256_in[1], zll_main_rotater256_in[0]};
  assign zll_main_rotater2529_in = {zll_main_rotater253_in[31], zll_main_rotater253_in[30], zll_main_rotater253_in[29], zll_main_rotater253_in[28], zll_main_rotater253_in[27], zll_main_rotater253_in[26], zll_main_rotater253_in[25], zll_main_rotater253_in[24], zll_main_rotater253_in[23], zll_main_rotater253_in[22], zll_main_rotater253_in[21], zll_main_rotater253_in[20], zll_main_rotater253_in[8], zll_main_rotater253_in[19], zll_main_rotater253_in[18], zll_main_rotater253_in[17], zll_main_rotater253_in[16], zll_main_rotater253_in[15], zll_main_rotater253_in[14], zll_main_rotater253_in[13], zll_main_rotater253_in[12], zll_main_rotater253_in[11], zll_main_rotater253_in[10], zll_main_rotater253_in[9], zll_main_rotater253_in[7], zll_main_rotater253_in[6], zll_main_rotater253_in[5], zll_main_rotater253_in[4], zll_main_rotater253_in[3], zll_main_rotater253_in[2], zll_main_rotater253_in[1], zll_main_rotater253_in[0]};
  assign zll_main_rotater2519_in = {zll_main_rotater2529_in[31], zll_main_rotater2529_in[30], zll_main_rotater2529_in[29], zll_main_rotater2529_in[28], zll_main_rotater2529_in[27], zll_main_rotater2529_in[26], zll_main_rotater2529_in[25], zll_main_rotater2529_in[24], zll_main_rotater2529_in[23], zll_main_rotater2529_in[22], zll_main_rotater2529_in[7], zll_main_rotater2529_in[21], zll_main_rotater2529_in[20], zll_main_rotater2529_in[19], zll_main_rotater2529_in[18], zll_main_rotater2529_in[17], zll_main_rotater2529_in[16], zll_main_rotater2529_in[15], zll_main_rotater2529_in[14], zll_main_rotater2529_in[13], zll_main_rotater2529_in[12], zll_main_rotater2529_in[11], zll_main_rotater2529_in[10], zll_main_rotater2529_in[9], zll_main_rotater2529_in[8], zll_main_rotater2529_in[6], zll_main_rotater2529_in[5], zll_main_rotater2529_in[4], zll_main_rotater2529_in[3], zll_main_rotater2529_in[2], zll_main_rotater2529_in[1], zll_main_rotater2529_in[0]};
  assign zll_main_rotater2514_in = {zll_main_rotater2519_in[31], zll_main_rotater2519_in[30], zll_main_rotater2519_in[29], zll_main_rotater2519_in[28], zll_main_rotater2519_in[27], zll_main_rotater2519_in[26], zll_main_rotater2519_in[25], zll_main_rotater2519_in[6], zll_main_rotater2519_in[24], zll_main_rotater2519_in[23], zll_main_rotater2519_in[22], zll_main_rotater2519_in[21], zll_main_rotater2519_in[20], zll_main_rotater2519_in[19], zll_main_rotater2519_in[18], zll_main_rotater2519_in[17], zll_main_rotater2519_in[16], zll_main_rotater2519_in[15], zll_main_rotater2519_in[14], zll_main_rotater2519_in[13], zll_main_rotater2519_in[12], zll_main_rotater2519_in[11], zll_main_rotater2519_in[10], zll_main_rotater2519_in[9], zll_main_rotater2519_in[8], zll_main_rotater2519_in[7], zll_main_rotater2519_in[5], zll_main_rotater2519_in[4], zll_main_rotater2519_in[3], zll_main_rotater2519_in[2], zll_main_rotater2519_in[1], zll_main_rotater2519_in[0]};
  assign zll_main_rotater2531_in = {zll_main_rotater2514_in[31], zll_main_rotater2514_in[30], zll_main_rotater2514_in[29], zll_main_rotater2514_in[28], zll_main_rotater2514_in[27], zll_main_rotater2514_in[26], zll_main_rotater2514_in[25], zll_main_rotater2514_in[24], zll_main_rotater2514_in[23], zll_main_rotater2514_in[22], zll_main_rotater2514_in[21], zll_main_rotater2514_in[20], zll_main_rotater2514_in[19], zll_main_rotater2514_in[18], zll_main_rotater2514_in[5], zll_main_rotater2514_in[17], zll_main_rotater2514_in[16], zll_main_rotater2514_in[15], zll_main_rotater2514_in[14], zll_main_rotater2514_in[13], zll_main_rotater2514_in[12], zll_main_rotater2514_in[11], zll_main_rotater2514_in[10], zll_main_rotater2514_in[9], zll_main_rotater2514_in[8], zll_main_rotater2514_in[7], zll_main_rotater2514_in[6], zll_main_rotater2514_in[4], zll_main_rotater2514_in[3], zll_main_rotater2514_in[2], zll_main_rotater2514_in[1], zll_main_rotater2514_in[0]};
  assign zll_main_rotater2517_in = {zll_main_rotater2531_in[31], zll_main_rotater2531_in[30], zll_main_rotater2531_in[29], zll_main_rotater2531_in[28], zll_main_rotater2531_in[27], zll_main_rotater2531_in[26], zll_main_rotater2531_in[25], zll_main_rotater2531_in[24], zll_main_rotater2531_in[23], zll_main_rotater2531_in[4], zll_main_rotater2531_in[22], zll_main_rotater2531_in[21], zll_main_rotater2531_in[20], zll_main_rotater2531_in[19], zll_main_rotater2531_in[18], zll_main_rotater2531_in[17], zll_main_rotater2531_in[16], zll_main_rotater2531_in[15], zll_main_rotater2531_in[14], zll_main_rotater2531_in[13], zll_main_rotater2531_in[12], zll_main_rotater2531_in[11], zll_main_rotater2531_in[10], zll_main_rotater2531_in[9], zll_main_rotater2531_in[8], zll_main_rotater2531_in[7], zll_main_rotater2531_in[6], zll_main_rotater2531_in[5], zll_main_rotater2531_in[3], zll_main_rotater2531_in[2], zll_main_rotater2531_in[1], zll_main_rotater2531_in[0]};
  assign zll_main_rotater2522_in = {zll_main_rotater2517_in[31], zll_main_rotater2517_in[30], zll_main_rotater2517_in[29], zll_main_rotater2517_in[28], zll_main_rotater2517_in[27], zll_main_rotater2517_in[26], zll_main_rotater2517_in[25], zll_main_rotater2517_in[24], zll_main_rotater2517_in[23], zll_main_rotater2517_in[22], zll_main_rotater2517_in[21], zll_main_rotater2517_in[20], zll_main_rotater2517_in[19], zll_main_rotater2517_in[18], zll_main_rotater2517_in[17], zll_main_rotater2517_in[16], zll_main_rotater2517_in[15], zll_main_rotater2517_in[14], zll_main_rotater2517_in[13], zll_main_rotater2517_in[3], zll_main_rotater2517_in[12], zll_main_rotater2517_in[11], zll_main_rotater2517_in[10], zll_main_rotater2517_in[9], zll_main_rotater2517_in[8], zll_main_rotater2517_in[7], zll_main_rotater2517_in[6], zll_main_rotater2517_in[5], zll_main_rotater2517_in[4], zll_main_rotater2517_in[2], zll_main_rotater2517_in[1], zll_main_rotater2517_in[0]};
  assign zll_main_rotater25_in = {zll_main_rotater2522_in[31], zll_main_rotater2522_in[30], zll_main_rotater2522_in[29], zll_main_rotater2522_in[28], zll_main_rotater2522_in[27], zll_main_rotater2522_in[26], zll_main_rotater2522_in[25], zll_main_rotater2522_in[24], zll_main_rotater2522_in[23], zll_main_rotater2522_in[22], zll_main_rotater2522_in[21], zll_main_rotater2522_in[20], zll_main_rotater2522_in[19], zll_main_rotater2522_in[18], zll_main_rotater2522_in[17], zll_main_rotater2522_in[16], zll_main_rotater2522_in[15], zll_main_rotater2522_in[14], zll_main_rotater2522_in[13], zll_main_rotater2522_in[12], zll_main_rotater2522_in[11], zll_main_rotater2522_in[10], zll_main_rotater2522_in[9], zll_main_rotater2522_in[8], zll_main_rotater2522_in[2], zll_main_rotater2522_in[7], zll_main_rotater2522_in[6], zll_main_rotater2522_in[5], zll_main_rotater2522_in[4], zll_main_rotater2522_in[3], zll_main_rotater2522_in[1], zll_main_rotater2522_in[0]};
  assign zll_main_rotater252_in = {zll_main_rotater25_in[31], zll_main_rotater25_in[30], zll_main_rotater25_in[29], zll_main_rotater25_in[28], zll_main_rotater25_in[27], zll_main_rotater25_in[26], zll_main_rotater25_in[25], zll_main_rotater25_in[24], zll_main_rotater25_in[23], zll_main_rotater25_in[22], zll_main_rotater25_in[21], zll_main_rotater25_in[20], zll_main_rotater25_in[19], zll_main_rotater25_in[18], zll_main_rotater25_in[17], zll_main_rotater25_in[16], zll_main_rotater25_in[1], zll_main_rotater25_in[15], zll_main_rotater25_in[14], zll_main_rotater25_in[13], zll_main_rotater25_in[12], zll_main_rotater25_in[11], zll_main_rotater25_in[10], zll_main_rotater25_in[9], zll_main_rotater25_in[8], zll_main_rotater25_in[7], zll_main_rotater25_in[6], zll_main_rotater25_in[5], zll_main_rotater25_in[4], zll_main_rotater25_in[3], zll_main_rotater25_in[2], zll_main_rotater25_in[0]};
  assign xorw32_inR1 = {extres, {zll_main_rotater252_in[17], zll_main_rotater252_in[20], zll_main_rotater252_in[8], zll_main_rotater252_in[28], zll_main_rotater252_in[4], zll_main_rotater252_in[29], zll_main_rotater252_in[13], zll_main_rotater252_in[9], zll_main_rotater252_in[1], zll_main_rotater252_in[27], zll_main_rotater252_in[21], zll_main_rotater252_in[5], zll_main_rotater252_in[31], zll_main_rotater252_in[2], zll_main_rotater252_in[3], zll_main_rotater252_in[18], zll_main_rotater252_in[14], zll_main_rotater252_in[19], zll_main_rotater252_in[24], zll_main_rotater252_in[16], zll_main_rotater252_in[22], zll_main_rotater252_in[11], zll_main_rotater252_in[6], zll_main_rotater252_in[15], zll_main_rotater252_in[0], zll_main_rotater252_in[30], zll_main_rotater252_in[25], zll_main_rotater252_in[7], zll_main_rotater252_in[23], zll_main_rotater252_in[12], zll_main_rotater252_in[26], zll_main_rotater252_in[10]}};
  xorW32  instR1 (xorw32_inR1[63:32], xorw32_inR1[31:0], extresR1[31:0]);
  assign res = extresR1;
endmodule

module ZLL_Main_dev32 (input logic [1029:0] arg0,
  output logic [1296:0] res);
  logic [1029:0] zll_main_dev54_in;
  logic [1029:0] zll_main_dev86_in;
  assign zll_main_dev54_in = arg0;
  assign zll_main_dev86_in = {zll_main_dev54_in[773:262], zll_main_dev54_in[1029:774], zll_main_dev54_in[261:6], zll_main_dev54_in[5:0]};
  assign res = {{10'h1, {9'h101{1'h0}}}, zll_main_dev86_in[517:262], zll_main_dev86_in[1029:518], zll_main_dev86_in[261:6], zll_main_dev86_in[5:0]};
endmodule

module Main_ch (input logic [31:0] arg0,
  input logic [31:0] arg1,
  input logic [31:0] arg2,
  output logic [31:0] res);
  logic [63:0] andw32_in;
  logic [31:0] extres;
  logic [31:0] notw32_in;
  logic [31:0] extresR1;
  logic [63:0] andw32_inR1;
  logic [31:0] extresR2;
  logic [63:0] xorw32_in;
  logic [31:0] extresR3;
  assign andw32_in = {arg0, arg1};
  andW32  inst (andw32_in[63:32], andw32_in[31:0], extres[31:0]);
  assign notw32_in = arg0;
  notW32  instR1 (notw32_in[31:0], extresR1[31:0]);
  assign andw32_inR1 = {extresR1, arg2};
  andW32  instR2 (andw32_inR1[63:32], andw32_inR1[31:0], extresR2[31:0]);
  assign xorw32_in = {extres, extresR2};
  xorW32  instR3 (xorw32_in[63:32], xorw32_in[31:0], extresR3[31:0]);
  assign res = extresR3;
endmodule